`default_nettype none
`timescale 1 ns / 1 ps

module rom(
    input  wire        clk,
    input  wire  [7:0] addr,
    output reg   [7:0] rddata
);

    always @(posedge clk) case (addr)
        8'h00: rddata <= 8'h3E;
        8'h01: rddata <= 8'h33;
        8'h02: rddata <= 8'hD3;
        8'h03: rddata <= 8'hF3;
        8'h04: rddata <= 8'h31;
        8'h05: rddata <= 8'h00;
        8'h06: rddata <= 8'h00;
        8'h07: rddata <= 8'hDB;
        8'h08: rddata <= 8'hFB;
        8'h09: rddata <= 8'hE6;
        8'h0A: rddata <= 8'h80;
        8'h0B: rddata <= 8'hF5;
        8'h0C: rddata <= 8'h3E;
        8'h0D: rddata <= 8'h06;
        8'h0E: rddata <= 8'hD3;
        8'h0F: rddata <= 8'hFB;
        8'h10: rddata <= 8'h3E;
        8'h11: rddata <= 8'h01;
        8'h12: rddata <= 8'hCD;
        8'h13: rddata <= 8'h6C;
        8'h14: rddata <= 8'h00;
        8'h15: rddata <= 8'h21;
        8'h16: rddata <= 8'h36;
        8'h17: rddata <= 8'h00;
        8'h18: rddata <= 8'hCD;
        8'h19: rddata <= 8'h4D;
        8'h1A: rddata <= 8'h00;
        8'h1B: rddata <= 8'h28;
        8'h1C: rddata <= 8'h06;
        8'h1D: rddata <= 8'h21;
        8'h1E: rddata <= 8'h40;
        8'h1F: rddata <= 8'h00;
        8'h20: rddata <= 8'hCD;
        8'h21: rddata <= 8'h4D;
        8'h22: rddata <= 8'h00;
        8'h23: rddata <= 8'h21;
        8'h24: rddata <= 8'h00;
        8'h25: rddata <= 8'hC0;
        8'h26: rddata <= 8'h11;
        8'h27: rddata <= 8'h00;
        8'h28: rddata <= 8'h30;
        8'h29: rddata <= 8'hCD;
        8'h2A: rddata <= 8'hA7;
        8'h2B: rddata <= 8'h00;
        8'h2C: rddata <= 8'hCD;
        8'h2D: rddata <= 8'h5F;
        8'h2E: rddata <= 8'h00;
        8'h2F: rddata <= 8'hE1;
        8'h30: rddata <= 8'hC3;
        8'h31: rddata <= 8'h00;
        8'h32: rddata <= 8'hC0;
        8'h33: rddata <= 8'hC3;
        8'h34: rddata <= 8'h33;
        8'h35: rddata <= 8'h00;
        8'h36: rddata <= 8'h2F;
        8'h37: rddata <= 8'h62;
        8'h38: rddata <= 8'h6F;
        8'h39: rddata <= 8'h6F;
        8'h3A: rddata <= 8'h74;
        8'h3B: rddata <= 8'h2E;
        8'h3C: rddata <= 8'h62;
        8'h3D: rddata <= 8'h69;
        8'h3E: rddata <= 8'h6E;
        8'h3F: rddata <= 8'h00;
        8'h40: rddata <= 8'h65;
        8'h41: rddata <= 8'h73;
        8'h42: rddata <= 8'h70;
        8'h43: rddata <= 8'h3A;
        8'h44: rddata <= 8'h62;
        8'h45: rddata <= 8'h6F;
        8'h46: rddata <= 8'h6F;
        8'h47: rddata <= 8'h74;
        8'h48: rddata <= 8'h2E;
        8'h49: rddata <= 8'h62;
        8'h4A: rddata <= 8'h69;
        8'h4B: rddata <= 8'h6E;
        8'h4C: rddata <= 8'h00;
        8'h4D: rddata <= 8'h3E;
        8'h4E: rddata <= 8'h10;
        8'h4F: rddata <= 8'hCD;
        8'h50: rddata <= 8'h6C;
        8'h51: rddata <= 8'h00;
        8'h52: rddata <= 8'h3E;
        8'h53: rddata <= 8'h00;
        8'h54: rddata <= 8'hCD;
        8'h55: rddata <= 8'h88;
        8'h56: rddata <= 8'h00;
        8'h57: rddata <= 8'hCD;
        8'h58: rddata <= 8'h9E;
        8'h59: rddata <= 8'h00;
        8'h5A: rddata <= 8'hCD;
        8'h5B: rddata <= 8'h7F;
        8'h5C: rddata <= 8'h00;
        8'h5D: rddata <= 8'hB7;
        8'h5E: rddata <= 8'hC9;
        8'h5F: rddata <= 8'h3E;
        8'h60: rddata <= 8'h11;
        8'h61: rddata <= 8'hCD;
        8'h62: rddata <= 8'h6C;
        8'h63: rddata <= 8'h00;
        8'h64: rddata <= 8'hAF;
        8'h65: rddata <= 8'hCD;
        8'h66: rddata <= 8'h88;
        8'h67: rddata <= 8'h00;
        8'h68: rddata <= 8'hCD;
        8'h69: rddata <= 8'h7F;
        8'h6A: rddata <= 8'h00;
        8'h6B: rddata <= 8'hC9;
        8'h6C: rddata <= 8'hF5;
        8'h6D: rddata <= 8'hDB;
        8'h6E: rddata <= 8'hF4;
        8'h6F: rddata <= 8'hE6;
        8'h70: rddata <= 8'h01;
        8'h71: rddata <= 8'h28;
        8'h72: rddata <= 8'h04;
        8'h73: rddata <= 8'hDB;
        8'h74: rddata <= 8'hF5;
        8'h75: rddata <= 8'h18;
        8'h76: rddata <= 8'hF6;
        8'h77: rddata <= 8'h3E;
        8'h78: rddata <= 8'h80;
        8'h79: rddata <= 8'hD3;
        8'h7A: rddata <= 8'hF4;
        8'h7B: rddata <= 8'hF1;
        8'h7C: rddata <= 8'hC3;
        8'h7D: rddata <= 8'h88;
        8'h7E: rddata <= 8'h00;
        8'h7F: rddata <= 8'hDB;
        8'h80: rddata <= 8'hF4;
        8'h81: rddata <= 8'hE6;
        8'h82: rddata <= 8'h01;
        8'h83: rddata <= 8'h28;
        8'h84: rddata <= 8'hFA;
        8'h85: rddata <= 8'hDB;
        8'h86: rddata <= 8'hF5;
        8'h87: rddata <= 8'hC9;
        8'h88: rddata <= 8'hF5;
        8'h89: rddata <= 8'hDB;
        8'h8A: rddata <= 8'hF4;
        8'h8B: rddata <= 8'hE6;
        8'h8C: rddata <= 8'h02;
        8'h8D: rddata <= 8'h20;
        8'h8E: rddata <= 8'hFA;
        8'h8F: rddata <= 8'hF1;
        8'h90: rddata <= 8'hD3;
        8'h91: rddata <= 8'hF5;
        8'h92: rddata <= 8'hC9;
        8'h93: rddata <= 8'h7A;
        8'h94: rddata <= 8'hB3;
        8'h95: rddata <= 8'hC8;
        8'h96: rddata <= 8'hCD;
        8'h97: rddata <= 8'h7F;
        8'h98: rddata <= 8'h00;
        8'h99: rddata <= 8'h77;
        8'h9A: rddata <= 8'h23;
        8'h9B: rddata <= 8'h1B;
        8'h9C: rddata <= 8'h18;
        8'h9D: rddata <= 8'hF5;
        8'h9E: rddata <= 8'h7E;
        8'h9F: rddata <= 8'h23;
        8'hA0: rddata <= 8'hCD;
        8'hA1: rddata <= 8'h88;
        8'hA2: rddata <= 8'h00;
        8'hA3: rddata <= 8'hB7;
        8'hA4: rddata <= 8'h20;
        8'hA5: rddata <= 8'hF8;
        8'hA6: rddata <= 8'hC9;
        8'hA7: rddata <= 8'h3E;
        8'hA8: rddata <= 8'h12;
        8'hA9: rddata <= 8'hCD;
        8'hAA: rddata <= 8'h6C;
        8'hAB: rddata <= 8'h00;
        8'hAC: rddata <= 8'hAF;
        8'hAD: rddata <= 8'hCD;
        8'hAE: rddata <= 8'h88;
        8'hAF: rddata <= 8'h00;
        8'hB0: rddata <= 8'h7B;
        8'hB1: rddata <= 8'hCD;
        8'hB2: rddata <= 8'h88;
        8'hB3: rddata <= 8'h00;
        8'hB4: rddata <= 8'h7A;
        8'hB5: rddata <= 8'hCD;
        8'hB6: rddata <= 8'h88;
        8'hB7: rddata <= 8'h00;
        8'hB8: rddata <= 8'hCD;
        8'hB9: rddata <= 8'h7F;
        8'hBA: rddata <= 8'h00;
        8'hBB: rddata <= 8'hB7;
        8'hBC: rddata <= 8'hC0;
        8'hBD: rddata <= 8'hCD;
        8'hBE: rddata <= 8'h7F;
        8'hBF: rddata <= 8'h00;
        8'hC0: rddata <= 8'h5F;
        8'hC1: rddata <= 8'hCD;
        8'hC2: rddata <= 8'h7F;
        8'hC3: rddata <= 8'h00;
        8'hC4: rddata <= 8'h57;
        8'hC5: rddata <= 8'hD5;
        8'hC6: rddata <= 8'h7A;
        8'hC7: rddata <= 8'hB3;
        8'hC8: rddata <= 8'h28;
        8'hC9: rddata <= 8'h08;
        8'hCA: rddata <= 8'hCD;
        8'hCB: rddata <= 8'h7F;
        8'hCC: rddata <= 8'h00;
        8'hCD: rddata <= 8'h77;
        8'hCE: rddata <= 8'h23;
        8'hCF: rddata <= 8'h1B;
        8'hD0: rddata <= 8'h18;
        8'hD1: rddata <= 8'hF4;
        8'hD2: rddata <= 8'hD1;
        8'hD3: rddata <= 8'hAF;
        8'hD4: rddata <= 8'hC9;
        default: rddata <= 8'h00;
    endcase

endmodule
