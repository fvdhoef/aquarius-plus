module colorram(
    input  wire       clk,

    input  wire [9:0] addr1,
    output reg  [7:0] rddata1,
    input  wire [7:0] wrdata1,
    input  wire       wren1,

    input  wire [9:0] addr2,
    output reg  [7:0] rddata2);

    reg [7:0] ram [1023:0];

    initial begin
        ram[   0] = 8'hDE; ram[   1] = 8'hE4; ram[   2] = 8'hE4; ram[   3] = 8'hE4;
        ram[   4] = 8'hE4; ram[   5] = 8'hE4; ram[   6] = 8'hE4; ram[   7] = 8'hE4;
        ram[   8] = 8'hE4; ram[   9] = 8'hE4; ram[  10] = 8'hE4; ram[  11] = 8'hE4;
        ram[  12] = 8'hE4; ram[  13] = 8'hE4; ram[  14] = 8'hE4; ram[  15] = 8'hE4;
        ram[  16] = 8'hE4; ram[  17] = 8'hE4; ram[  18] = 8'hE4; ram[  19] = 8'hE4;
        ram[  20] = 8'hE4; ram[  21] = 8'hE4; ram[  22] = 8'hE4; ram[  23] = 8'hE4;
        ram[  24] = 8'hE4; ram[  25] = 8'hE4; ram[  26] = 8'hE4; ram[  27] = 8'hE4;
        ram[  28] = 8'hE4; ram[  29] = 8'hE4; ram[  30] = 8'hE4; ram[  31] = 8'hE4;
        ram[  32] = 8'hE4; ram[  33] = 8'hE4; ram[  34] = 8'hE4; ram[  35] = 8'hE4;
        ram[  36] = 8'hE4; ram[  37] = 8'hE4; ram[  38] = 8'hE4; ram[  39] = 8'hE4;
        ram[  40] = 8'hE4; ram[  41] = 8'hE4; ram[  42] = 8'hE4; ram[  43] = 8'hE4;
        ram[  44] = 8'hE4; ram[  45] = 8'hE4; ram[  46] = 8'hE4; ram[  47] = 8'hE4;
        ram[  48] = 8'hE4; ram[  49] = 8'hE4; ram[  50] = 8'hE4; ram[  51] = 8'hE4;
        ram[  52] = 8'hE4; ram[  53] = 8'hE4; ram[  54] = 8'hE4; ram[  55] = 8'hE4;
        ram[  56] = 8'hE4; ram[  57] = 8'hE4; ram[  58] = 8'hE4; ram[  59] = 8'hE4;
        ram[  60] = 8'hE4; ram[  61] = 8'h74; ram[  62] = 8'hE4; ram[  63] = 8'hE4;
        ram[  64] = 8'hE4; ram[  65] = 8'h74; ram[  66] = 8'h84; ram[  67] = 8'h74;
        ram[  68] = 8'h74; ram[  69] = 8'hE4; ram[  70] = 8'hE4; ram[  71] = 8'hE4;
        ram[  72] = 8'hE4; ram[  73] = 8'hE4; ram[  74] = 8'hE4; ram[  75] = 8'hE4;
        ram[  76] = 8'hE4; ram[  77] = 8'h74; ram[  78] = 8'hE4; ram[  79] = 8'hE4;
        ram[  80] = 8'hE4; ram[  81] = 8'h74; ram[  82] = 8'hE4; ram[  83] = 8'hE4;
        ram[  84] = 8'hE4; ram[  85] = 8'hE4; ram[  86] = 8'hE4; ram[  87] = 8'h74;
        ram[  88] = 8'hE4; ram[  89] = 8'hE4; ram[  90] = 8'hE4; ram[  91] = 8'hE4;
        ram[  92] = 8'h74; ram[  93] = 8'hE4; ram[  94] = 8'hE4; ram[  95] = 8'hE4;
        ram[  96] = 8'hE4; ram[  97] = 8'hE4; ram[  98] = 8'h74; ram[  99] = 8'hE4;
        ram[ 100] = 8'hE4; ram[ 101] = 8'hE4; ram[ 102] = 8'hE4; ram[ 103] = 8'hE4;
        ram[ 104] = 8'hE4; ram[ 105] = 8'h0E; ram[ 106] = 8'hE0; ram[ 107] = 8'hEE;
        ram[ 108] = 8'hEE; ram[ 109] = 8'hE4; ram[ 110] = 8'hE4; ram[ 111] = 8'h74;
        ram[ 112] = 8'hE4; ram[ 113] = 8'hE4; ram[ 114] = 8'hE4; ram[ 115] = 8'hE4;
        ram[ 116] = 8'hE4; ram[ 117] = 8'hE4; ram[ 118] = 8'hE4; ram[ 119] = 8'h74;
        ram[ 120] = 8'hE4; ram[ 121] = 8'hE4; ram[ 122] = 8'hE4; ram[ 123] = 8'h34;
        ram[ 124] = 8'h34; ram[ 125] = 8'hE4; ram[ 126] = 8'hE4; ram[ 127] = 8'hE4;
        ram[ 128] = 8'hE4; ram[ 129] = 8'hE4; ram[ 130] = 8'hE4; ram[ 131] = 8'hE4;
        ram[ 132] = 8'hE4; ram[ 133] = 8'hE4; ram[ 134] = 8'h04; ram[ 135] = 8'h04;
        ram[ 136] = 8'h04; ram[ 137] = 8'h04; ram[ 138] = 8'h04; ram[ 139] = 8'h04;
        ram[ 140] = 8'h04; ram[ 141] = 8'h04; ram[ 142] = 8'h04; ram[ 143] = 8'h04;
        ram[ 144] = 8'hE4; ram[ 145] = 8'h0E; ram[ 146] = 8'hE0; ram[ 147] = 8'hEE;
        ram[ 148] = 8'hEE; ram[ 149] = 8'hE4; ram[ 150] = 8'hE4; ram[ 151] = 8'hE4;
        ram[ 152] = 8'hE4; ram[ 153] = 8'hE4; ram[ 154] = 8'hE4; ram[ 155] = 8'hE4;
        ram[ 156] = 8'hE4; ram[ 157] = 8'hE4; ram[ 158] = 8'hE4; ram[ 159] = 8'hE4;
        ram[ 160] = 8'hE4; ram[ 161] = 8'hE4; ram[ 162] = 8'h34; ram[ 163] = 8'hC4;
        ram[ 164] = 8'hC4; ram[ 165] = 8'h34; ram[ 166] = 8'hE4; ram[ 167] = 8'hE4;
        ram[ 168] = 8'hE4; ram[ 169] = 8'hE4; ram[ 170] = 8'hE4; ram[ 171] = 8'hE4;
        ram[ 172] = 8'h74; ram[ 173] = 8'h87; ram[ 174] = 8'h87; ram[ 175] = 8'h87;
        ram[ 176] = 8'h87; ram[ 177] = 8'h87; ram[ 178] = 8'h87; ram[ 179] = 8'h87;
        ram[ 180] = 8'h87; ram[ 181] = 8'h87; ram[ 182] = 8'h87; ram[ 183] = 8'h87;
        ram[ 184] = 8'h87; ram[ 185] = 8'h0E; ram[ 186] = 8'hE0; ram[ 187] = 8'hEE;
        ram[ 188] = 8'h7E; ram[ 189] = 8'h87; ram[ 190] = 8'h87; ram[ 191] = 8'h87;
        ram[ 192] = 8'hE7; ram[ 193] = 8'hE4; ram[ 194] = 8'hE4; ram[ 195] = 8'hE4;
        ram[ 196] = 8'h74; ram[ 197] = 8'hE4; ram[ 198] = 8'hE4; ram[ 199] = 8'hE4;
        ram[ 200] = 8'hE4; ram[ 201] = 8'hE4; ram[ 202] = 8'h34; ram[ 203] = 8'hC4;
        ram[ 204] = 8'hC4; ram[ 205] = 8'h34; ram[ 206] = 8'hE4; ram[ 207] = 8'h74;
        ram[ 208] = 8'hE4; ram[ 209] = 8'hE4; ram[ 210] = 8'hE4; ram[ 211] = 8'h74;
        ram[ 212] = 8'h87; ram[ 213] = 8'h87; ram[ 214] = 8'h7F; ram[ 215] = 8'h87;
        ram[ 216] = 8'h7F; ram[ 217] = 8'h7F; ram[ 218] = 8'h7F; ram[ 219] = 8'h7F;
        ram[ 220] = 8'h7F; ram[ 221] = 8'h87; ram[ 222] = 8'h7F; ram[ 223] = 8'h7F;
        ram[ 224] = 8'h7F; ram[ 225] = 8'h0E; ram[ 226] = 8'hE0; ram[ 227] = 8'h7E;
        ram[ 228] = 8'h7F; ram[ 229] = 8'h7F; ram[ 230] = 8'h7F; ram[ 231] = 8'hE7;
        ram[ 232] = 8'hEF; ram[ 233] = 8'hEF; ram[ 234] = 8'hE4; ram[ 235] = 8'hE4;
        ram[ 236] = 8'hE4; ram[ 237] = 8'hE4; ram[ 238] = 8'hE4; ram[ 239] = 8'hE4;
        ram[ 240] = 8'hE4; ram[ 241] = 8'hE4; ram[ 242] = 8'hE4; ram[ 243] = 8'h34;
        ram[ 244] = 8'h34; ram[ 245] = 8'hE4; ram[ 246] = 8'hE4; ram[ 247] = 8'hE4;
        ram[ 248] = 8'hE4; ram[ 249] = 8'hE4; ram[ 250] = 8'h74; ram[ 251] = 8'h87;
        ram[ 252] = 8'h87; ram[ 253] = 8'h7F; ram[ 254] = 8'h7F; ram[ 255] = 8'h7F;
        ram[ 256] = 8'h87; ram[ 257] = 8'h7F; ram[ 258] = 8'h87; ram[ 259] = 8'h7F;
        ram[ 260] = 8'h7F; ram[ 261] = 8'h7F; ram[ 262] = 8'h7F; ram[ 263] = 8'h87;
        ram[ 264] = 8'h7F; ram[ 265] = 8'h7F; ram[ 266] = 8'h7F; ram[ 267] = 8'h87;
        ram[ 268] = 8'h7F; ram[ 269] = 8'h7F; ram[ 270] = 8'hE7; ram[ 271] = 8'hEF;
        ram[ 272] = 8'hF0; ram[ 273] = 8'hF0; ram[ 274] = 8'hEF; ram[ 275] = 8'hE4;
        ram[ 276] = 8'hE4; ram[ 277] = 8'h74; ram[ 278] = 8'hE4; ram[ 279] = 8'h74;
        ram[ 280] = 8'hE4; ram[ 281] = 8'hE4; ram[ 282] = 8'hE4; ram[ 283] = 8'hE4;
        ram[ 284] = 8'hE4; ram[ 285] = 8'hE4; ram[ 286] = 8'hE4; ram[ 287] = 8'hE4;
        ram[ 288] = 8'hE4; ram[ 289] = 8'h74; ram[ 290] = 8'h87; ram[ 291] = 8'h87;
        ram[ 292] = 8'h7F; ram[ 293] = 8'h7F; ram[ 294] = 8'h87; ram[ 295] = 8'h7F;
        ram[ 296] = 8'h7F; ram[ 297] = 8'h7F; ram[ 298] = 8'h7F; ram[ 299] = 8'h87;
        ram[ 300] = 8'h7F; ram[ 301] = 8'h7F; ram[ 302] = 8'h87; ram[ 303] = 8'h7F;
        ram[ 304] = 8'h7F; ram[ 305] = 8'h87; ram[ 306] = 8'h7F; ram[ 307] = 8'h7F;
        ram[ 308] = 8'h7F; ram[ 309] = 8'hE7; ram[ 310] = 8'hEF; ram[ 311] = 8'hEF;
        ram[ 312] = 8'h0F; ram[ 313] = 8'h0F; ram[ 314] = 8'hEF; ram[ 315] = 8'hEF;
        ram[ 316] = 8'hE4; ram[ 317] = 8'hE4; ram[ 318] = 8'hE4; ram[ 319] = 8'hE4;
        ram[ 320] = 8'hE4; ram[ 321] = 8'hE4; ram[ 322] = 8'hE4; ram[ 323] = 8'hE4;
        ram[ 324] = 8'h74; ram[ 325] = 8'hE4; ram[ 326] = 8'hE4; ram[ 327] = 8'hE4;
        ram[ 328] = 8'h74; ram[ 329] = 8'h87; ram[ 330] = 8'h87; ram[ 331] = 8'h7F;
        ram[ 332] = 8'h7F; ram[ 333] = 8'h87; ram[ 334] = 8'h87; ram[ 335] = 8'h7F;
        ram[ 336] = 8'h7F; ram[ 337] = 8'h7F; ram[ 338] = 8'h7F; ram[ 339] = 8'h7F;
        ram[ 340] = 8'h7F; ram[ 341] = 8'h7F; ram[ 342] = 8'h7F; ram[ 343] = 8'h7F;
        ram[ 344] = 8'h7F; ram[ 345] = 8'h7F; ram[ 346] = 8'h7F; ram[ 347] = 8'h7F;
        ram[ 348] = 8'hE7; ram[ 349] = 8'hEF; ram[ 350] = 8'hEF; ram[ 351] = 8'hEF;
        ram[ 352] = 8'hEF; ram[ 353] = 8'hEF; ram[ 354] = 8'hEF; ram[ 355] = 8'hEF;
        ram[ 356] = 8'hEF; ram[ 357] = 8'hE4; ram[ 358] = 8'hE4; ram[ 359] = 8'hE4;
        ram[ 360] = 8'hE4; ram[ 361] = 8'hE4; ram[ 362] = 8'hE4; ram[ 363] = 8'hE4;
        ram[ 364] = 8'hE4; ram[ 365] = 8'hE4; ram[ 366] = 8'hE4; ram[ 367] = 8'hE4;
        ram[ 368] = 8'h0E; ram[ 369] = 8'hE0; ram[ 370] = 8'hE0; ram[ 371] = 8'hE0;
        ram[ 372] = 8'h7E; ram[ 373] = 8'h7E; ram[ 374] = 8'hE0; ram[ 375] = 8'hE0;
        ram[ 376] = 8'h7E; ram[ 377] = 8'hE0; ram[ 378] = 8'hE7; ram[ 379] = 8'h7F;
        ram[ 380] = 8'hE7; ram[ 381] = 8'hE0; ram[ 382] = 8'hE0; ram[ 383] = 8'hE0;
        ram[ 384] = 8'h7E; ram[ 385] = 8'h7E; ram[ 386] = 8'h7E; ram[ 387] = 8'hE0;
        ram[ 388] = 8'h0E; ram[ 389] = 8'hEF; ram[ 390] = 8'h7E; ram[ 391] = 8'h7E;
        ram[ 392] = 8'hEF; ram[ 393] = 8'h7E; ram[ 394] = 8'h7E; ram[ 395] = 8'h7E;
        ram[ 396] = 8'h7E; ram[ 397] = 8'hEB; ram[ 398] = 8'hE4; ram[ 399] = 8'hE4;
        ram[ 400] = 8'h74; ram[ 401] = 8'hE4; ram[ 402] = 8'hE4; ram[ 403] = 8'h14;
        ram[ 404] = 8'hE4; ram[ 405] = 8'hE4; ram[ 406] = 8'hE4; ram[ 407] = 8'hE4;
        ram[ 408] = 8'h0E; ram[ 409] = 8'hEF; ram[ 410] = 8'hEF; ram[ 411] = 8'hEF;
        ram[ 412] = 8'hEF; ram[ 413] = 8'h0E; ram[ 414] = 8'h0E; ram[ 415] = 8'h0E;
        ram[ 416] = 8'hEF; ram[ 417] = 8'hEF; ram[ 418] = 8'hEF; ram[ 419] = 8'h7E;
        ram[ 420] = 8'hEF; ram[ 421] = 8'hEF; ram[ 422] = 8'hEF; ram[ 423] = 8'h0E;
        ram[ 424] = 8'h0E; ram[ 425] = 8'h0E; ram[ 426] = 8'hEF; ram[ 427] = 8'hEF;
        ram[ 428] = 8'h0E; ram[ 429] = 8'hEF; ram[ 430] = 8'hEF; ram[ 431] = 8'h0E;
        ram[ 432] = 8'h0E; ram[ 433] = 8'h0E; ram[ 434] = 8'h0E; ram[ 435] = 8'h0E;
        ram[ 436] = 8'hEF; ram[ 437] = 8'hE0; ram[ 438] = 8'hE4; ram[ 439] = 8'h74;
        ram[ 440] = 8'hE4; ram[ 441] = 8'hE4; ram[ 442] = 8'hE4; ram[ 443] = 8'h34;
        ram[ 444] = 8'hE4; ram[ 445] = 8'hE4; ram[ 446] = 8'hE4; ram[ 447] = 8'hE4;
        ram[ 448] = 8'h0E; ram[ 449] = 8'hEF; ram[ 450] = 8'hEF; ram[ 451] = 8'hEF;
        ram[ 452] = 8'hE0; ram[ 453] = 8'hC7; ram[ 454] = 8'hC7; ram[ 455] = 8'hC7;
        ram[ 456] = 8'h0E; ram[ 457] = 8'hEF; ram[ 458] = 8'hEF; ram[ 459] = 8'h1E;
        ram[ 460] = 8'hEF; ram[ 461] = 8'hEF; ram[ 462] = 8'hE0; ram[ 463] = 8'hC7;
        ram[ 464] = 8'hC7; ram[ 465] = 8'hC7; ram[ 466] = 8'h0E; ram[ 467] = 8'hEF;
        ram[ 468] = 8'h0E; ram[ 469] = 8'hEF; ram[ 470] = 8'hE0; ram[ 471] = 8'h0C;
        ram[ 472] = 8'h7C; ram[ 473] = 8'h0C; ram[ 474] = 8'h7C; ram[ 475] = 8'h0C;
        ram[ 476] = 8'h0E; ram[ 477] = 8'hE0; ram[ 478] = 8'hE4; ram[ 479] = 8'hE4;
        ram[ 480] = 8'hE4; ram[ 481] = 8'hE4; ram[ 482] = 8'h24; ram[ 483] = 8'h12;
        ram[ 484] = 8'h24; ram[ 485] = 8'hE4; ram[ 486] = 8'hE4; ram[ 487] = 8'hE4;
        ram[ 488] = 8'h0E; ram[ 489] = 8'hEF; ram[ 490] = 8'hEF; ram[ 491] = 8'hEF;
        ram[ 492] = 8'hE0; ram[ 493] = 8'h7C; ram[ 494] = 8'h7C; ram[ 495] = 8'h7C;
        ram[ 496] = 8'h0E; ram[ 497] = 8'hEF; ram[ 498] = 8'h1E; ram[ 499] = 8'hDE;
        ram[ 500] = 8'h1E; ram[ 501] = 8'hEF; ram[ 502] = 8'hE0; ram[ 503] = 8'h7C;
        ram[ 504] = 8'h7C; ram[ 505] = 8'h7C; ram[ 506] = 8'h0E; ram[ 507] = 8'hEF;
        ram[ 508] = 8'h0E; ram[ 509] = 8'hEF; ram[ 510] = 8'hE0; ram[ 511] = 8'h7C;
        ram[ 512] = 8'h0C; ram[ 513] = 8'h0C; ram[ 514] = 8'h0C; ram[ 515] = 8'h7C;
        ram[ 516] = 8'h0E; ram[ 517] = 8'hE0; ram[ 518] = 8'hE4; ram[ 519] = 8'hE4;
        ram[ 520] = 8'hE4; ram[ 521] = 8'h24; ram[ 522] = 8'h12; ram[ 523] = 8'h22;
        ram[ 524] = 8'h42; ram[ 525] = 8'h24; ram[ 526] = 8'hE4; ram[ 527] = 8'hE4;
        ram[ 528] = 8'h0E; ram[ 529] = 8'hEF; ram[ 530] = 8'hEF; ram[ 531] = 8'hEF;
        ram[ 532] = 8'hE0; ram[ 533] = 8'h5C; ram[ 534] = 8'h5C; ram[ 535] = 8'hDC;
        ram[ 536] = 8'h0E; ram[ 537] = 8'hEF; ram[ 538] = 8'hE0; ram[ 539] = 8'hE0;
        ram[ 540] = 8'hE0; ram[ 541] = 8'hEF; ram[ 542] = 8'hE0; ram[ 543] = 8'h1C;
        ram[ 544] = 8'h4C; ram[ 545] = 8'h7C; ram[ 546] = 8'h0E; ram[ 547] = 8'hEF;
        ram[ 548] = 8'h0E; ram[ 549] = 8'hEF; ram[ 550] = 8'hE0; ram[ 551] = 8'h7C;
        ram[ 552] = 8'h0C; ram[ 553] = 8'h0C; ram[ 554] = 8'h0C; ram[ 555] = 8'h7C;
        ram[ 556] = 8'h0E; ram[ 557] = 8'hE0; ram[ 558] = 8'h74; ram[ 559] = 8'hE4;
        ram[ 560] = 8'hE4; ram[ 561] = 8'h24; ram[ 562] = 8'h72; ram[ 563] = 8'h12;
        ram[ 564] = 8'h24; ram[ 565] = 8'h24; ram[ 566] = 8'hE4; ram[ 567] = 8'h74;
        ram[ 568] = 8'h0E; ram[ 569] = 8'hEF; ram[ 570] = 8'hEF; ram[ 571] = 8'hEF;
        ram[ 572] = 8'hEF; ram[ 573] = 8'hE0; ram[ 574] = 8'hE0; ram[ 575] = 8'hE0;
        ram[ 576] = 8'hEF; ram[ 577] = 8'hE0; ram[ 578] = 8'hC7; ram[ 579] = 8'h7C;
        ram[ 580] = 8'hC7; ram[ 581] = 8'h0E; ram[ 582] = 8'hEF; ram[ 583] = 8'hE0;
        ram[ 584] = 8'hE0; ram[ 585] = 8'hE0; ram[ 586] = 8'hEF; ram[ 587] = 8'hEF;
        ram[ 588] = 8'h0E; ram[ 589] = 8'hEF; ram[ 590] = 8'hEF; ram[ 591] = 8'hE0;
        ram[ 592] = 8'hE0; ram[ 593] = 8'hE0; ram[ 594] = 8'hE0; ram[ 595] = 8'hE0;
        ram[ 596] = 8'h6E; ram[ 597] = 8'h6E; ram[ 598] = 8'h64; ram[ 599] = 8'hE4;
        ram[ 600] = 8'hE4; ram[ 601] = 8'h24; ram[ 602] = 8'h22; ram[ 603] = 8'h22;
        ram[ 604] = 8'h52; ram[ 605] = 8'h24; ram[ 606] = 8'hE4; ram[ 607] = 8'hE4;
        ram[ 608] = 8'h0E; ram[ 609] = 8'hEF; ram[ 610] = 8'hEF; ram[ 611] = 8'hEF;
        ram[ 612] = 8'hEF; ram[ 613] = 8'hEF; ram[ 614] = 8'hEF; ram[ 615] = 8'hEF;
        ram[ 616] = 8'hEF; ram[ 617] = 8'hE0; ram[ 618] = 8'h7C; ram[ 619] = 8'h1C;
        ram[ 620] = 8'h7C; ram[ 621] = 8'h0E; ram[ 622] = 8'hEF; ram[ 623] = 8'hEF;
        ram[ 624] = 8'hEF; ram[ 625] = 8'hEF; ram[ 626] = 8'hEF; ram[ 627] = 8'hEF;
        ram[ 628] = 8'h0E; ram[ 629] = 8'h7E; ram[ 630] = 8'h7E; ram[ 631] = 8'hEF;
        ram[ 632] = 8'hEF; ram[ 633] = 8'hEF; ram[ 634] = 8'hEF; ram[ 635] = 8'hEF;
        ram[ 636] = 8'hEF; ram[ 637] = 8'h7E; ram[ 638] = 8'hE4; ram[ 639] = 8'hE4;
        ram[ 640] = 8'hE4; ram[ 641] = 8'h24; ram[ 642] = 8'h42; ram[ 643] = 8'h32;
        ram[ 644] = 8'h24; ram[ 645] = 8'h24; ram[ 646] = 8'hE4; ram[ 647] = 8'hE4;
        ram[ 648] = 8'h0E; ram[ 649] = 8'hEF; ram[ 650] = 8'hEF; ram[ 651] = 8'h7E;
        ram[ 652] = 8'h7E; ram[ 653] = 8'hEF; ram[ 654] = 8'hEF; ram[ 655] = 8'hEF;
        ram[ 656] = 8'hEF; ram[ 657] = 8'hE0; ram[ 658] = 8'h7C; ram[ 659] = 8'h1C;
        ram[ 660] = 8'h7C; ram[ 661] = 8'h0E; ram[ 662] = 8'hEF; ram[ 663] = 8'hEF;
        ram[ 664] = 8'hEF; ram[ 665] = 8'hEF; ram[ 666] = 8'hEF; ram[ 667] = 8'h7E;
        ram[ 668] = 8'h07; ram[ 669] = 8'h07; ram[ 670] = 8'h07; ram[ 671] = 8'h7E;
        ram[ 672] = 8'hEF; ram[ 673] = 8'hEF; ram[ 674] = 8'hEF; ram[ 675] = 8'hEF;
        ram[ 676] = 8'h7E; ram[ 677] = 8'hD7; ram[ 678] = 8'h74; ram[ 679] = 8'hE4;
        ram[ 680] = 8'h74; ram[ 681] = 8'hE4; ram[ 682] = 8'hE4; ram[ 683] = 8'hE4;
        ram[ 684] = 8'hE4; ram[ 685] = 8'hE4; ram[ 686] = 8'hE4; ram[ 687] = 8'h74;
        ram[ 688] = 8'h0E; ram[ 689] = 8'h7E; ram[ 690] = 8'h7E; ram[ 691] = 8'h07;
        ram[ 692] = 8'h07; ram[ 693] = 8'h7E; ram[ 694] = 8'h7E; ram[ 695] = 8'h7E;
        ram[ 696] = 8'hEF; ram[ 697] = 8'hE0; ram[ 698] = 8'h7C; ram[ 699] = 8'hFC;
        ram[ 700] = 8'h7C; ram[ 701] = 8'h0E; ram[ 702] = 8'hEF; ram[ 703] = 8'hEF;
        ram[ 704] = 8'h7E; ram[ 705] = 8'hEF; ram[ 706] = 8'h7E; ram[ 707] = 8'h07;
        ram[ 708] = 8'h07; ram[ 709] = 8'h87; ram[ 710] = 8'h07; ram[ 711] = 8'h07;
        ram[ 712] = 8'h7E; ram[ 713] = 8'h7E; ram[ 714] = 8'hEF; ram[ 715] = 8'hEF;
        ram[ 716] = 8'h7E; ram[ 717] = 8'h07; ram[ 718] = 8'h74; ram[ 719] = 8'hE4;
        ram[ 720] = 8'h87; ram[ 721] = 8'h07; ram[ 722] = 8'h07; ram[ 723] = 8'h87;
        ram[ 724] = 8'h07; ram[ 725] = 8'h07; ram[ 726] = 8'h07; ram[ 727] = 8'h07;
        ram[ 728] = 8'h07; ram[ 729] = 8'h07; ram[ 730] = 8'h07; ram[ 731] = 8'h87;
        ram[ 732] = 8'h07; ram[ 733] = 8'h07; ram[ 734] = 8'h07; ram[ 735] = 8'h07;
        ram[ 736] = 8'h87; ram[ 737] = 8'h8F; ram[ 738] = 8'h08; ram[ 739] = 8'h8F;
        ram[ 740] = 8'h8F; ram[ 741] = 8'h8F; ram[ 742] = 8'h78; ram[ 743] = 8'h07;
        ram[ 744] = 8'h07; ram[ 745] = 8'h07; ram[ 746] = 8'h07; ram[ 747] = 8'h07;
        ram[ 748] = 8'h07; ram[ 749] = 8'h07; ram[ 750] = 8'h07; ram[ 751] = 8'h07;
        ram[ 752] = 8'h07; ram[ 753] = 8'h07; ram[ 754] = 8'h07; ram[ 755] = 8'h07;
        ram[ 756] = 8'h07; ram[ 757] = 8'h07; ram[ 758] = 8'h07; ram[ 759] = 8'h07;
        ram[ 760] = 8'h07; ram[ 761] = 8'h87; ram[ 762] = 8'h87; ram[ 763] = 8'h07;
        ram[ 764] = 8'h07; ram[ 765] = 8'h07; ram[ 766] = 8'h87; ram[ 767] = 8'h07;
        ram[ 768] = 8'h07; ram[ 769] = 8'h87; ram[ 770] = 8'h87; ram[ 771] = 8'h07;
        ram[ 772] = 8'h07; ram[ 773] = 8'h87; ram[ 774] = 8'h07; ram[ 775] = 8'h87;
        ram[ 776] = 8'h8F; ram[ 777] = 8'h08; ram[ 778] = 8'h08; ram[ 779] = 8'h8F;
        ram[ 780] = 8'h8F; ram[ 781] = 8'h78; ram[ 782] = 8'h07; ram[ 783] = 8'h87;
        ram[ 784] = 8'h07; ram[ 785] = 8'h87; ram[ 786] = 8'h07; ram[ 787] = 8'h87;
        ram[ 788] = 8'h07; ram[ 789] = 8'h87; ram[ 790] = 8'h07; ram[ 791] = 8'h07;
        ram[ 792] = 8'h87; ram[ 793] = 8'h07; ram[ 794] = 8'h87; ram[ 795] = 8'h07;
        ram[ 796] = 8'h87; ram[ 797] = 8'h07; ram[ 798] = 8'h07; ram[ 799] = 8'h87;
        ram[ 800] = 8'h07; ram[ 801] = 8'h07; ram[ 802] = 8'h87; ram[ 803] = 8'h07;
        ram[ 804] = 8'h07; ram[ 805] = 8'h87; ram[ 806] = 8'h07; ram[ 807] = 8'h87;
        ram[ 808] = 8'h07; ram[ 809] = 8'h07; ram[ 810] = 8'h07; ram[ 811] = 8'h07;
        ram[ 812] = 8'h87; ram[ 813] = 8'h07; ram[ 814] = 8'h87; ram[ 815] = 8'h08;
        ram[ 816] = 8'h08; ram[ 817] = 8'h08; ram[ 818] = 8'h08; ram[ 819] = 8'h8F;
        ram[ 820] = 8'h78; ram[ 821] = 8'h07; ram[ 822] = 8'h07; ram[ 823] = 8'h07;
        ram[ 824] = 8'h07; ram[ 825] = 8'h07; ram[ 826] = 8'h87; ram[ 827] = 8'h07;
        ram[ 828] = 8'h07; ram[ 829] = 8'h07; ram[ 830] = 8'h87; ram[ 831] = 8'h07;
        ram[ 832] = 8'h87; ram[ 833] = 8'h07; ram[ 834] = 8'h07; ram[ 835] = 8'h87;
        ram[ 836] = 8'h07; ram[ 837] = 8'h07; ram[ 838] = 8'h07; ram[ 839] = 8'h07;
        ram[ 840] = 8'h87; ram[ 841] = 8'h07; ram[ 842] = 8'h07; ram[ 843] = 8'h07;
        ram[ 844] = 8'h07; ram[ 845] = 8'h07; ram[ 846] = 8'h87; ram[ 847] = 8'h07;
        ram[ 848] = 8'h07; ram[ 849] = 8'h07; ram[ 850] = 8'h87; ram[ 851] = 8'h07;
        ram[ 852] = 8'h07; ram[ 853] = 8'h87; ram[ 854] = 8'h8F; ram[ 855] = 8'h08;
        ram[ 856] = 8'h08; ram[ 857] = 8'h08; ram[ 858] = 8'h8F; ram[ 859] = 8'h78;
        ram[ 860] = 8'h07; ram[ 861] = 8'h87; ram[ 862] = 8'h07; ram[ 863] = 8'h87;
        ram[ 864] = 8'h07; ram[ 865] = 8'h07; ram[ 866] = 8'h07; ram[ 867] = 8'h07;
        ram[ 868] = 8'h07; ram[ 869] = 8'h07; ram[ 870] = 8'h07; ram[ 871] = 8'h87;
        ram[ 872] = 8'h07; ram[ 873] = 8'h07; ram[ 874] = 8'h07; ram[ 875] = 8'h07;
        ram[ 876] = 8'h07; ram[ 877] = 8'h07; ram[ 878] = 8'h87; ram[ 879] = 8'h07;
        ram[ 880] = 8'h8F; ram[ 881] = 8'h8F; ram[ 882] = 8'h8F; ram[ 883] = 8'h8F;
        ram[ 884] = 8'h8F; ram[ 885] = 8'h8F; ram[ 886] = 8'h8F; ram[ 887] = 8'h8F;
        ram[ 888] = 8'h8F; ram[ 889] = 8'h8F; ram[ 890] = 8'h8F; ram[ 891] = 8'h8F;
        ram[ 892] = 8'h8F; ram[ 893] = 8'h58; ram[ 894] = 8'h08; ram[ 895] = 8'h08;
        ram[ 896] = 8'h08; ram[ 897] = 8'h28; ram[ 898] = 8'h8F; ram[ 899] = 8'h8F;
        ram[ 900] = 8'h8F; ram[ 901] = 8'h8F; ram[ 902] = 8'h8F; ram[ 903] = 8'h8F;
        ram[ 904] = 8'h8F; ram[ 905] = 8'h8F; ram[ 906] = 8'h8F; ram[ 907] = 8'h8F;
        ram[ 908] = 8'h8F; ram[ 909] = 8'h8F; ram[ 910] = 8'h8F; ram[ 911] = 8'h8F;
        ram[ 912] = 8'h8F; ram[ 913] = 8'h8F; ram[ 914] = 8'h8F; ram[ 915] = 8'h8F;
        ram[ 916] = 8'h8F; ram[ 917] = 8'h8F; ram[ 918] = 8'h8F; ram[ 919] = 8'h8F;
        ram[ 920] = 8'h48; ram[ 921] = 8'h08; ram[ 922] = 8'h38; ram[ 923] = 8'h08;
        ram[ 924] = 8'h08; ram[ 925] = 8'h38; ram[ 926] = 8'h08; ram[ 927] = 8'h08;
        ram[ 928] = 8'h38; ram[ 929] = 8'h08; ram[ 930] = 8'h08; ram[ 931] = 8'h38;
        ram[ 932] = 8'h08; ram[ 933] = 8'h08; ram[ 934] = 8'h38; ram[ 935] = 8'h08;
        ram[ 936] = 8'h08; ram[ 937] = 8'hD8; ram[ 938] = 8'h08; ram[ 939] = 8'h08;
        ram[ 940] = 8'h38; ram[ 941] = 8'h08; ram[ 942] = 8'h08; ram[ 943] = 8'h38;
        ram[ 944] = 8'h08; ram[ 945] = 8'h08; ram[ 946] = 8'h38; ram[ 947] = 8'hD8;
        ram[ 948] = 8'h08; ram[ 949] = 8'h38; ram[ 950] = 8'h08; ram[ 951] = 8'h08;
        ram[ 952] = 8'h38; ram[ 953] = 8'h08; ram[ 954] = 8'h08; ram[ 955] = 8'h38;
        ram[ 956] = 8'h08; ram[ 957] = 8'h08; ram[ 958] = 8'h38; ram[ 959] = 8'h08;
        ram[ 960] = 8'h08; ram[ 961] = 8'h08; ram[ 962] = 8'h08; ram[ 963] = 8'h08;
        ram[ 964] = 8'h08; ram[ 965] = 8'h08; ram[ 966] = 8'h08; ram[ 967] = 8'hD8;
        ram[ 968] = 8'h08; ram[ 969] = 8'h08; ram[ 970] = 8'h08; ram[ 971] = 8'h08;
        ram[ 972] = 8'h08; ram[ 973] = 8'h08; ram[ 974] = 8'h08; ram[ 975] = 8'h08;
        ram[ 976] = 8'h08; ram[ 977] = 8'h08; ram[ 978] = 8'h08; ram[ 979] = 8'h08;
        ram[ 980] = 8'h08; ram[ 981] = 8'h18; ram[ 982] = 8'h08; ram[ 983] = 8'h08;
        ram[ 984] = 8'h08; ram[ 985] = 8'h08; ram[ 986] = 8'h08; ram[ 987] = 8'h08;
        ram[ 988] = 8'h08; ram[ 989] = 8'h08; ram[ 990] = 8'h08; ram[ 991] = 8'h08;
        ram[ 992] = 8'h08; ram[ 993] = 8'h08; ram[ 994] = 8'h08; ram[ 995] = 8'h08;
        ram[ 996] = 8'h48; ram[ 997] = 8'h08; ram[ 998] = 8'h08; ram[ 999] = 8'h08;
        ram[1000] = 8'h00; ram[1001] = 8'h00; ram[1002] = 8'h00; ram[1003] = 8'h00;
        ram[1004] = 8'h00; ram[1005] = 8'h00; ram[1006] = 8'h00; ram[1007] = 8'h00;
        ram[1008] = 8'h00; ram[1009] = 8'h00; ram[1010] = 8'h00; ram[1011] = 8'h00;
        ram[1012] = 8'h00; ram[1013] = 8'h00; ram[1014] = 8'h00; ram[1015] = 8'h00;
        ram[1016] = 8'h00; ram[1017] = 8'h00; ram[1018] = 8'h00; ram[1019] = 8'h00;
        ram[1020] = 8'h00; ram[1021] = 8'h00; ram[1022] = 8'h00; ram[1023] = 8'h00;
    end

    always @(posedge clk)
    begin
        if (wren1) ram[addr1] = wrdata1;
        rddata1 <= ram[addr1];
    end

    always @(posedge clk)
    begin
        rddata2 <= ram[addr2];
    end

endmodule
