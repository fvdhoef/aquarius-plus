`default_nettype none
`timescale 1 ns / 1 ps

module charram(
    input  wire        clk1,
    input  wire [10:0] addr1,
    output wire  [7:0] rddata1,
    input  wire  [7:0] wrdata1,
    input  wire        wren1,

    input  wire        clk2,
    input  wire [10:0] addr2,
    output wire  [7:0] rddata2);

    wire [0:0] dopa, dopb;  // unused

    RAMB16_S9_S9 #(
        .INIT_A(9'h000),                // Value of output RAM registers on Port A at startup
        .INIT_B(9'h000),                // Value of output RAM registers on Port B at startup
        .SRVAL_A(9'h000),               // Port A output value upon SSR assertion
        .SRVAL_B(9'h000),               // Port B output value upon SSR assertion
        .WRITE_MODE_A("WRITE_FIRST"),   // WRITE_FIRST, READ_FIRST or NO_CHANGE
        .WRITE_MODE_B("WRITE_FIRST"),   // WRITE_FIRST, READ_FIRST or NO_CHANGE
        .SIM_COLLISION_CHECK("NONE"),   // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL"

        // The following INIT_xx declarations specify the initial contents of the RAM
        .INIT_00(256'h00041C542C50286400041C542C504844001C08442C50484400AC60207820203C),
        .INIT_01(256'h002040FFFF402000000402FFFF0204003C4299A1A199423C000010007C001000),
        .INIT_02(256'hF0E0F0B81C0E0400002070381D0F070F183C5A181818181818181818185A3C18),
        .INIT_03(256'h30303030303CFCFCFFFFFF7E003C3C0000040E1CB8F0E0F00F070F1D38702000),
        .INIT_04(256'hDBBDFF7E003C3C003C3C3C3C3C3C3C3C0C0C0C0C0C3C3F3F0000003C3C3C3CFF),
        .INIT_05(256'hDCDF7939003C38003838181C1E1B3E7C7F7C7838003C3800C3C3C3E766663C7E),
        .INIT_06(256'h000000000F0F0F0F0F0F0F0F00000000DB99BDE724663C180080C3F33B1F3F7C),
        .INIT_07(256'hFFFFFFFF000000000F0F0F0FF0F0F0F000000000F0F0F0F0F0F0F0F000000000),
        .INIT_08(256'h0028287C287C2828000000000028282800100010101010100000000000000000),
        .INIT_09(256'h00000000001008080034485420505020000C4C20100864600010781438503C10),
        .INIT_0A(256'h000010107C101000001054381038541000100804040408100010204040402010),
        .INIT_0B(256'h00004020100804000010000000000000000000007C0000000020101000000000),
        .INIT_0C(256'h003844041808047C007C402018044438003810101010301000384464544C4438),
        .INIT_0D(256'h002020201008047C003844447840201C003844040478407C0008087C48281808),
        .INIT_0E(256'h00201010001000000000001000100000007008043C4444380038444438444438),
        .INIT_0F(256'h001000101008443800201008040810200000007C007C00000008102040201008),
        .INIT_10(256'h003844404040443800784444784444780044447C44442810003C40585C544438),
        .INIT_11(256'h003C444C4040403C004040407840407C007C40407840407C0078444444444478),
        .INIT_12(256'h004448506050484400384404040404040038101010101038004444447C444444),
        .INIT_13(256'h00384444444444380044444C546444440044444454546C44007C404040404040),
        .INIT_14(256'h0038440438404438004448507844447800344854444444380040404078444478),
        .INIT_15(256'h00446C545444444400102844444444440038444444444444001010101010107C),
        .INIT_16(256'h007C60606060607C007C40201008047C00101010102844440044442810284444),
        .INIT_17(256'h007C0000000000000000004428100000007C0C0C0C0C0C7C0000040810204000),
        .INIT_18(256'h001C2020201C0000005864446458404000344C444C3400000000000000102020),
        .INIT_19(256'h38043C444C34000000101010381010080038407C4438000000344C444C340404),
        .INIT_1A(256'h0044487050484040300808080808000800381010103000100044444444784040),
        .INIT_1B(256'h0038444444380000004444444478000000525252526C00000038101010101030),
        .INIT_1C(256'h00780438403C0000004040406058000006344C444C3400004058644464580000),
        .INIT_1D(256'h002C5252525200000010282844440000003C44444444000000101010107C1010),
        .INIT_1E(256'h000C10102010100C007C2010087C000038043C24242400000044281028440000),
        .INIT_1F(256'hFFFFFFFFFFFFFFFF000000403804000000601010081010600010101000101010),
        .INIT_20(256'h1C1C183878D87C3EFE3E1E1C003C1C008080808080808080FFFFFFFFFFFFFF00),
        .INIT_21(256'h00183C7E7E3C180055AA55AA55AA55AA50A050A050A050A055AA55AA00000000),
        .INIT_22(256'h18183C7EFFDB183C3C18DBFF7E3C1818FFFFFFFFFFFF0000FFFF000000000000),
        .INIT_23(256'hFFFF7E7E3C3C1818C0F0FCFFFFFCF0C00001C3CFDCF8FC3E3BFB9E9C003C1C00),
        .INIT_24(256'hBCBCFF3D013C4A3C3D3DFFBC803C523CFEFEFEFEFEFEFEFEFF00000000000000),
        .INIT_25(256'hC0C0C0C0C0C0C0C03C7EFFFFFFFF7E3C050A050A050A050A0000000055AA55AA),
        .INIT_26(256'h0C1C39FFFF391C0C30389CFFFF9C3830F8F8F8F8F8F8F8F8E0E0E0E0E0E0E0E0),
        .INIT_27(256'h18183C3C7E7EFFFF030F3FFFFF3F0F0300667E42C3FF18000018FFC3427E6600),
        .INIT_28(256'h0000000000FFFFFF00000000000F0F0F0000000000F0F0F00000000000000000),
        .INIT_29(256'h000000F0F0FFFFFF000000F0F00F0F0F000000F0F0F0F0F0000000F0F0000000),
        .INIT_2A(256'h0000000F0FFFFFFF0000000F0F0F0F0F0000000F0FF0F0F00000000F0F000000),
        .INIT_2B(256'h000000FFFFFFFFFF000000FFFF0F0F0F000000FFFFF0F0F0000000FFFF000000),
        .INIT_2C(256'hF0F0F00000FFFFFFF0F0F000000F0F0FF0F0F00000F0F0F0F0F0F00000000000),
        .INIT_2D(256'hF0F0F0F0F0FFFFFFF0F0F0F0F00F0F0FF0F0F0F0F0F0F0F0F0F0F0F0F0000000),
        .INIT_2E(256'hF0F0F00F0FFFFFFFF0F0F00F0F0F0F0FF0F0F00F0FF0F0F0F0F0F00F0F000000),
        .INIT_2F(256'hF0F0F0FFFFFFFFFFF0F0F0FFFF0F0F0FF0F0F0FFFFF0F0F0F0F0F0FFFF000000),
        .INIT_30(256'hFCFCFCFCFCFCFCFC000000003C7EFFFFFFFEFCF8F0E0C080FF7F3F1F0F070301),
        .INIT_31(256'h0000000003070F0F0000001818000000183C7EFFFF7E3C1800003C3C3C3C0000),
        .INIT_32(256'h03070F0F0F0F07038040201008040201F0F0E0C000000000181818FFFF181818),
        .INIT_33(256'h0000001F1F181818181818F8F80000001818181F1F181818000000FFFF181818),
        .INIT_34(256'h0004345C3A2C1000FFFF7E3C000000004A23B411C42D44520208401180042009),
        .INIT_35(256'h0F0F07030000000018181818181818183C1842E742183C1818183C7EFFFFFF66),
        .INIT_36(256'hC0E0F0F0F0F0E0C0010204081020408000000000C0E0F0F08142241818244281),
        .INIT_37(256'h000000F8F81818181818181F1F000000181818F8F8181818181818FFFF000000),
        .INIT_38(256'h0F0F0F0000FFFFFF0F0F0F00000F0F0F0F0F0F0000F0F0F00F0F0F0000000000),
        .INIT_39(256'h0F0F0FF0F0FFFFFF0F0F0FF0F00F0F0F0F0F0FF0F0F0F0F00F0F0FF0F0000000),
        .INIT_3A(256'h0F0F0F0F0FFFFFFF0F0F0F0F0F0F0F0F0F0F0F0F0FF0F0F00F0F0F0F0F000000),
        .INIT_3B(256'h0F0F0FFFFFFFFFFF0F0F0FFFFF0F0F0F0F0F0FFFFFF0F0F00F0F0FFFFF000000),
        .INIT_3C(256'hFFFFFF0000FFFFFFFFFFFF00000F0F0FFFFFFF0000F0F0F0FFFFFF0000000000),
        .INIT_3D(256'hFFFFFFF0F0FFFFFFFFFFFFF0F00F0F0FFFFFFFF0F0F0F0F0FFFFFFF0F0000000),
        .INIT_3E(256'hFFFFFF0F0FFFFFFFFFFFFF0F0F0F0F0FFFFFFF0F0FF0F0F0FFFFFF0F0F000000),
        .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0F0F0FFFFFFFFFFFF0F0F0FFFFFFFFFF000000)
    )
    
    RAMB16_S9_S9_inst(
        .CLKA(clk1),
        .SSRA(1'b0),
        .ADDRA(addr1),
        .DOA(rddata1),
        .DOPA(dopa),
        .DIA(wrdata1),
        .DIPA(1'b0),
        .ENA(1'b1),
        .WEA(wren1),

        .CLKB(clk2),
        .SSRB(1'b0),
        .ADDRB(addr2),
        .DOB(rddata2),
        .DOPB(dopb),
        .DIB(8'b0),
        .DIPB(1'b0),
        .ENB(1'b1),
        .WEB(1'b0)
    );

endmodule
