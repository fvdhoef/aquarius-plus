`default_nettype none
`timescale 1 ns / 1 ps

module rom(
    input  wire        clk,
    input  wire [12:0] addr,
    output reg   [7:0] rddata
);

    always @(posedge clk) case (addr)
        13'h00: rddata <= 8'hF3;
        13'h01: rddata <= 8'hED;
        13'h02: rddata <= 8'h56;
        13'h03: rddata <= 8'h31;
        13'h04: rddata <= 8'h00;
        13'h05: rddata <= 8'hDF;
        13'h06: rddata <= 8'h21;
        13'h07: rddata <= 8'h00;
        13'h08: rddata <= 8'hC0;
        13'h09: rddata <= 8'h11;
        13'h0A: rddata <= 8'h01;
        13'h0B: rddata <= 8'hC0;
        13'h0C: rddata <= 8'h01;
        13'h0D: rddata <= 8'hFF;
        13'h0E: rddata <= 8'h1F;
        13'h0F: rddata <= 8'h36;
        13'h10: rddata <= 8'h00;
        13'h11: rddata <= 8'hED;
        13'h12: rddata <= 8'hB0;
        13'h13: rddata <= 8'hAF;
        13'h14: rddata <= 8'h32;
        13'h15: rddata <= 8'hFD;
        13'h16: rddata <= 8'hFF;
        13'h17: rddata <= 8'h3E;
        13'h18: rddata <= 8'h01;
        13'h19: rddata <= 8'hCD;
        13'h1A: rddata <= 8'hF7;
        13'h1B: rddata <= 8'h0F;
        13'h1C: rddata <= 8'hC3;
        13'h1D: rddata <= 8'h1F;
        13'h1E: rddata <= 8'h00;
        13'h1F: rddata <= 8'hCD;
        13'h20: rddata <= 8'h09;
        13'h21: rddata <= 8'h03;
        13'h22: rddata <= 8'hCD;
        13'h23: rddata <= 8'h86;
        13'h24: rddata <= 8'h0F;
        13'h25: rddata <= 8'hCD;
        13'h26: rddata <= 8'hFB;
        13'h27: rddata <= 8'h00;
        13'h28: rddata <= 8'hCD;
        13'h29: rddata <= 8'h2D;
        13'h2A: rddata <= 8'h01;
        13'h2B: rddata <= 8'hCD;
        13'h2C: rddata <= 8'h7A;
        13'h2D: rddata <= 8'h0F;
        13'h2E: rddata <= 8'hCD;
        13'h2F: rddata <= 8'h86;
        13'h30: rddata <= 8'h0F;
        13'h31: rddata <= 8'hCD;
        13'h32: rddata <= 8'hFB;
        13'h33: rddata <= 8'h00;
        13'h34: rddata <= 8'hC3;
        13'h35: rddata <= 8'h66;
        13'h36: rddata <= 8'h00;
        13'h37: rddata <= 8'hCD;
        13'h38: rddata <= 8'h32;
        13'h39: rddata <= 8'h10;
        13'h3A: rddata <= 8'hCD;
        13'h3B: rddata <= 8'h3A;
        13'h3C: rddata <= 8'h10;
        13'h3D: rddata <= 8'h3A;
        13'h3E: rddata <= 8'h02;
        13'h3F: rddata <= 8'hC0;
        13'h40: rddata <= 8'h47;
        13'h41: rddata <= 8'h04;
        13'h42: rddata <= 8'h05;
        13'h43: rddata <= 8'h28;
        13'h44: rddata <= 8'h07;
        13'h45: rddata <= 8'h0E;
        13'h46: rddata <= 8'h16;
        13'h47: rddata <= 8'hCD;
        13'h48: rddata <= 8'h5A;
        13'h49: rddata <= 8'h00;
        13'h4A: rddata <= 8'h18;
        13'h4B: rddata <= 8'hF6;
        13'h4C: rddata <= 8'h3A;
        13'h4D: rddata <= 8'h03;
        13'h4E: rddata <= 8'hC0;
        13'h4F: rddata <= 8'h4F;
        13'h50: rddata <= 8'hCD;
        13'h51: rddata <= 8'h5A;
        13'h52: rddata <= 8'h00;
        13'h53: rddata <= 8'hCD;
        13'h54: rddata <= 8'h46;
        13'h55: rddata <= 8'h10;
        13'h56: rddata <= 8'hCD;
        13'h57: rddata <= 8'h32;
        13'h58: rddata <= 8'h10;
        13'h59: rddata <= 8'hC9;
        13'h5A: rddata <= 8'h79;
        13'h5B: rddata <= 8'hB7;
        13'h5C: rddata <= 8'hC8;
        13'h5D: rddata <= 8'hC5;
        13'h5E: rddata <= 8'hCD;
        13'h5F: rddata <= 8'h46;
        13'h60: rddata <= 8'h10;
        13'h61: rddata <= 8'hC1;
        13'h62: rddata <= 8'h0D;
        13'h63: rddata <= 8'hC8;
        13'h64: rddata <= 8'h18;
        13'h65: rddata <= 8'hF7;
        13'h66: rddata <= 8'hCD;
        13'h67: rddata <= 8'h37;
        13'h68: rddata <= 8'h00;
        13'h69: rddata <= 8'hAF;
        13'h6A: rddata <= 8'h32;
        13'h6B: rddata <= 8'h00;
        13'h6C: rddata <= 8'hC0;
        13'h6D: rddata <= 8'h3E;
        13'h6E: rddata <= 8'h08;
        13'h6F: rddata <= 8'h32;
        13'h70: rddata <= 8'h01;
        13'h71: rddata <= 8'hC0;
        13'h72: rddata <= 8'hCD;
        13'h73: rddata <= 8'h9D;
        13'h74: rddata <= 8'h0F;
        13'h75: rddata <= 8'h21;
        13'h76: rddata <= 8'h92;
        13'h77: rddata <= 8'h00;
        13'h78: rddata <= 8'hCD;
        13'h79: rddata <= 8'hEE;
        13'h7A: rddata <= 8'h0F;
        13'h7B: rddata <= 8'hCD;
        13'h7C: rddata <= 8'hD3;
        13'h7D: rddata <= 8'h02;
        13'h7E: rddata <= 8'hCD;
        13'h7F: rddata <= 8'h9D;
        13'h80: rddata <= 8'h00;
        13'h81: rddata <= 8'hCD;
        13'h82: rddata <= 8'h32;
        13'h83: rddata <= 8'h10;
        13'h84: rddata <= 8'h11;
        13'h85: rddata <= 8'h00;
        13'h86: rddata <= 8'hD0;
        13'h87: rddata <= 8'h21;
        13'h88: rddata <= 8'hD3;
        13'h89: rddata <= 8'h10;
        13'h8A: rddata <= 8'h01;
        13'h8B: rddata <= 8'h13;
        13'h8C: rddata <= 8'h00;
        13'h8D: rddata <= 8'hED;
        13'h8E: rddata <= 8'hB0;
        13'h8F: rddata <= 8'hC3;
        13'h90: rddata <= 8'h00;
        13'h91: rddata <= 8'hD0;
        13'h92: rddata <= 8'h4C;
        13'h93: rddata <= 8'h6F;
        13'h94: rddata <= 8'h61;
        13'h95: rddata <= 8'h64;
        13'h96: rddata <= 8'h69;
        13'h97: rddata <= 8'h6E;
        13'h98: rddata <= 8'h67;
        13'h99: rddata <= 8'h3A;
        13'h9A: rddata <= 8'h0A;
        13'h9B: rddata <= 8'h0A;
        13'h9C: rddata <= 8'h00;
        13'h9D: rddata <= 8'hCD;
        13'h9E: rddata <= 8'h32;
        13'h9F: rddata <= 8'h10;
        13'hA0: rddata <= 8'h3E;
        13'hA1: rddata <= 8'h10;
        13'hA2: rddata <= 8'hCD;
        13'hA3: rddata <= 8'hF7;
        13'hA4: rddata <= 8'h0F;
        13'hA5: rddata <= 8'h3E;
        13'hA6: rddata <= 8'h00;
        13'hA7: rddata <= 8'hCD;
        13'hA8: rddata <= 8'h13;
        13'hA9: rddata <= 8'h10;
        13'hAA: rddata <= 8'h21;
        13'hAB: rddata <= 8'h12;
        13'hAC: rddata <= 8'hC0;
        13'hAD: rddata <= 8'h7E;
        13'hAE: rddata <= 8'h23;
        13'hAF: rddata <= 8'hCD;
        13'hB0: rddata <= 8'h13;
        13'hB1: rddata <= 8'h10;
        13'hB2: rddata <= 8'hB7;
        13'hB3: rddata <= 8'h20;
        13'hB4: rddata <= 8'hF8;
        13'hB5: rddata <= 8'hCD;
        13'hB6: rddata <= 8'h0A;
        13'hB7: rddata <= 8'h10;
        13'hB8: rddata <= 8'h3A;
        13'hB9: rddata <= 8'h0F;
        13'hBA: rddata <= 8'hC0;
        13'hBB: rddata <= 8'hCB;
        13'hBC: rddata <= 8'h4F;
        13'hBD: rddata <= 8'h28;
        13'hBE: rddata <= 8'h1B;
        13'hBF: rddata <= 8'h3E;
        13'hC0: rddata <= 8'h14;
        13'hC1: rddata <= 8'hCD;
        13'hC2: rddata <= 8'hF7;
        13'hC3: rddata <= 8'h0F;
        13'hC4: rddata <= 8'hAF;
        13'hC5: rddata <= 8'hCD;
        13'hC6: rddata <= 8'h13;
        13'hC7: rddata <= 8'h10;
        13'hC8: rddata <= 8'hCD;
        13'hC9: rddata <= 8'h13;
        13'hCA: rddata <= 8'h10;
        13'hCB: rddata <= 8'h3E;
        13'hCC: rddata <= 8'h02;
        13'hCD: rddata <= 8'hCD;
        13'hCE: rddata <= 8'h13;
        13'hCF: rddata <= 8'h10;
        13'hD0: rddata <= 8'hAF;
        13'hD1: rddata <= 8'hCD;
        13'hD2: rddata <= 8'h13;
        13'hD3: rddata <= 8'h10;
        13'hD4: rddata <= 8'hCD;
        13'hD5: rddata <= 8'h13;
        13'hD6: rddata <= 8'h10;
        13'hD7: rddata <= 8'hCD;
        13'hD8: rddata <= 8'h0A;
        13'hD9: rddata <= 8'h10;
        13'hDA: rddata <= 8'hAF;
        13'hDB: rddata <= 8'h32;
        13'hDC: rddata <= 8'hFE;
        13'hDD: rddata <= 8'hFF;
        13'hDE: rddata <= 8'h21;
        13'hDF: rddata <= 8'h00;
        13'hE0: rddata <= 8'h40;
        13'hE1: rddata <= 8'h11;
        13'hE2: rddata <= 8'h00;
        13'hE3: rddata <= 8'h40;
        13'hE4: rddata <= 8'hCD;
        13'hE5: rddata <= 8'hA8;
        13'hE6: rddata <= 8'h10;
        13'hE7: rddata <= 8'h7A;
        13'hE8: rddata <= 8'hFE;
        13'hE9: rddata <= 8'h40;
        13'hEA: rddata <= 8'h20;
        13'hEB: rddata <= 8'h0E;
        13'hEC: rddata <= 8'h3E;
        13'hED: rddata <= 8'h2E;
        13'hEE: rddata <= 8'hCD;
        13'hEF: rddata <= 8'hB6;
        13'hF0: rddata <= 8'h0F;
        13'hF1: rddata <= 8'h3A;
        13'hF2: rddata <= 8'hFE;
        13'hF3: rddata <= 8'hFF;
        13'hF4: rddata <= 8'h3C;
        13'hF5: rddata <= 8'h32;
        13'hF6: rddata <= 8'hFE;
        13'hF7: rddata <= 8'hFF;
        13'hF8: rddata <= 8'h18;
        13'hF9: rddata <= 8'hE4;
        13'hFA: rddata <= 8'hC9;
        13'hFB: rddata <= 8'hAF;
        13'hFC: rddata <= 8'h32;
        13'hFD: rddata <= 8'h00;
        13'hFE: rddata <= 8'hC0;
        13'hFF: rddata <= 8'h32;
        13'h100: rddata <= 8'h01;
        13'h101: rddata <= 8'hC0;
        13'h102: rddata <= 8'hCD;
        13'h103: rddata <= 8'h9D;
        13'h104: rddata <= 8'h0F;
        13'h105: rddata <= 8'h21;
        13'h106: rddata <= 8'h0C;
        13'h107: rddata <= 8'h01;
        13'h108: rddata <= 8'hCD;
        13'h109: rddata <= 8'hEE;
        13'h10A: rddata <= 8'h0F;
        13'h10B: rddata <= 8'hC9;
        13'h10C: rddata <= 8'h3C;
        13'h10D: rddata <= 8'h3C;
        13'h10E: rddata <= 8'h3C;
        13'h10F: rddata <= 8'h3C;
        13'h110: rddata <= 8'h20;
        13'h111: rddata <= 8'h41;
        13'h112: rddata <= 8'h71;
        13'h113: rddata <= 8'h75;
        13'h114: rddata <= 8'h61;
        13'h115: rddata <= 8'h72;
        13'h116: rddata <= 8'h69;
        13'h117: rddata <= 8'h75;
        13'h118: rddata <= 8'h73;
        13'h119: rddata <= 8'h20;
        13'h11A: rddata <= 8'h4D;
        13'h11B: rddata <= 8'h61;
        13'h11C: rddata <= 8'h73;
        13'h11D: rddata <= 8'h74;
        13'h11E: rddata <= 8'h65;
        13'h11F: rddata <= 8'h72;
        13'h120: rddata <= 8'h20;
        13'h121: rddata <= 8'h53;
        13'h122: rddata <= 8'h79;
        13'h123: rddata <= 8'h73;
        13'h124: rddata <= 8'h74;
        13'h125: rddata <= 8'h65;
        13'h126: rddata <= 8'h6D;
        13'h127: rddata <= 8'h20;
        13'h128: rddata <= 8'h3E;
        13'h129: rddata <= 8'h3E;
        13'h12A: rddata <= 8'h3E;
        13'h12B: rddata <= 8'h3E;
        13'h12C: rddata <= 8'h00;
        13'h12D: rddata <= 8'hCD;
        13'h12E: rddata <= 8'h27;
        13'h12F: rddata <= 8'h02;
        13'h130: rddata <= 8'hCD;
        13'h131: rddata <= 8'h14;
        13'h132: rddata <= 8'h02;
        13'h133: rddata <= 8'h3A;
        13'h134: rddata <= 8'h05;
        13'h135: rddata <= 8'hC0;
        13'h136: rddata <= 8'hCB;
        13'h137: rddata <= 8'h5F;
        13'h138: rddata <= 8'h20;
        13'h139: rddata <= 8'h16;
        13'h13A: rddata <= 8'hCB;
        13'h13B: rddata <= 8'h57;
        13'h13C: rddata <= 8'h20;
        13'h13D: rddata <= 8'h17;
        13'h13E: rddata <= 8'hCB;
        13'h13F: rddata <= 8'h47;
        13'h140: rddata <= 8'h20;
        13'h141: rddata <= 8'h18;
        13'h142: rddata <= 8'hCB;
        13'h143: rddata <= 8'h4F;
        13'h144: rddata <= 8'h20;
        13'h145: rddata <= 8'h19;
        13'h146: rddata <= 8'hCB;
        13'h147: rddata <= 8'h67;
        13'h148: rddata <= 8'h20;
        13'h149: rddata <= 8'h1A;
        13'h14A: rddata <= 8'hCB;
        13'h14B: rddata <= 8'h6F;
        13'h14C: rddata <= 8'h20;
        13'h14D: rddata <= 8'h1B;
        13'h14E: rddata <= 8'h18;
        13'h14F: rddata <= 8'hE0;
        13'h150: rddata <= 8'hCD;
        13'h151: rddata <= 8'h03;
        13'h152: rddata <= 8'h02;
        13'h153: rddata <= 8'h18;
        13'h154: rddata <= 8'hDB;
        13'h155: rddata <= 8'hCD;
        13'h156: rddata <= 8'hF3;
        13'h157: rddata <= 8'h01;
        13'h158: rddata <= 8'h18;
        13'h159: rddata <= 8'hD6;
        13'h15A: rddata <= 8'hCD;
        13'h15B: rddata <= 8'hBA;
        13'h15C: rddata <= 8'h01;
        13'h15D: rddata <= 8'h18;
        13'h15E: rddata <= 8'hD1;
        13'h15F: rddata <= 8'hCD;
        13'h160: rddata <= 8'hD3;
        13'h161: rddata <= 8'h01;
        13'h162: rddata <= 8'h18;
        13'h163: rddata <= 8'hCC;
        13'h164: rddata <= 8'hCD;
        13'h165: rddata <= 8'h9B;
        13'h166: rddata <= 8'h01;
        13'h167: rddata <= 8'h18;
        13'h168: rddata <= 8'hC7;
        13'h169: rddata <= 8'h3A;
        13'h16A: rddata <= 8'h07;
        13'h16B: rddata <= 8'hC0;
        13'h16C: rddata <= 8'hB7;
        13'h16D: rddata <= 8'h28;
        13'h16E: rddata <= 8'hC1;
        13'h16F: rddata <= 8'hCD;
        13'h170: rddata <= 8'h37;
        13'h171: rddata <= 8'h00;
        13'h172: rddata <= 8'h3A;
        13'h173: rddata <= 8'h0D;
        13'h174: rddata <= 8'hC0;
        13'h175: rddata <= 8'hCB;
        13'h176: rddata <= 8'h47;
        13'h177: rddata <= 8'hC8;
        13'h178: rddata <= 8'hCD;
        13'h179: rddata <= 8'h7D;
        13'h17A: rddata <= 8'h01;
        13'h17B: rddata <= 8'h18;
        13'h17C: rddata <= 8'hB3;
        13'h17D: rddata <= 8'h3E;
        13'h17E: rddata <= 8'h1C;
        13'h17F: rddata <= 8'hCD;
        13'h180: rddata <= 8'hF7;
        13'h181: rddata <= 8'h0F;
        13'h182: rddata <= 8'h21;
        13'h183: rddata <= 8'h12;
        13'h184: rddata <= 8'hC0;
        13'h185: rddata <= 8'h7E;
        13'h186: rddata <= 8'h23;
        13'h187: rddata <= 8'hCD;
        13'h188: rddata <= 8'h13;
        13'h189: rddata <= 8'h10;
        13'h18A: rddata <= 8'hB7;
        13'h18B: rddata <= 8'h20;
        13'h18C: rddata <= 8'hF8;
        13'h18D: rddata <= 8'hCD;
        13'h18E: rddata <= 8'h0A;
        13'h18F: rddata <= 8'h10;
        13'h190: rddata <= 8'hAF;
        13'h191: rddata <= 8'h32;
        13'h192: rddata <= 8'h02;
        13'h193: rddata <= 8'hC0;
        13'h194: rddata <= 8'h32;
        13'h195: rddata <= 8'h03;
        13'h196: rddata <= 8'hC0;
        13'h197: rddata <= 8'hCD;
        13'h198: rddata <= 8'h27;
        13'h199: rddata <= 8'h02;
        13'h19A: rddata <= 8'hC9;
        13'h19B: rddata <= 8'h3E;
        13'h19C: rddata <= 8'h1C;
        13'h19D: rddata <= 8'hCD;
        13'h19E: rddata <= 8'hF7;
        13'h19F: rddata <= 8'h0F;
        13'h1A0: rddata <= 8'h3E;
        13'h1A1: rddata <= 8'h2E;
        13'h1A2: rddata <= 8'hCD;
        13'h1A3: rddata <= 8'h13;
        13'h1A4: rddata <= 8'h10;
        13'h1A5: rddata <= 8'hCD;
        13'h1A6: rddata <= 8'h13;
        13'h1A7: rddata <= 8'h10;
        13'h1A8: rddata <= 8'hAF;
        13'h1A9: rddata <= 8'hCD;
        13'h1AA: rddata <= 8'h13;
        13'h1AB: rddata <= 8'h10;
        13'h1AC: rddata <= 8'hCD;
        13'h1AD: rddata <= 8'h0A;
        13'h1AE: rddata <= 8'h10;
        13'h1AF: rddata <= 8'hAF;
        13'h1B0: rddata <= 8'h32;
        13'h1B1: rddata <= 8'h02;
        13'h1B2: rddata <= 8'hC0;
        13'h1B3: rddata <= 8'h32;
        13'h1B4: rddata <= 8'h03;
        13'h1B5: rddata <= 8'hC0;
        13'h1B6: rddata <= 8'hCD;
        13'h1B7: rddata <= 8'h27;
        13'h1B8: rddata <= 8'h02;
        13'h1B9: rddata <= 8'hC9;
        13'h1BA: rddata <= 8'h3A;
        13'h1BB: rddata <= 8'h03;
        13'h1BC: rddata <= 8'hC0;
        13'h1BD: rddata <= 8'hB7;
        13'h1BE: rddata <= 8'h28;
        13'h1BF: rddata <= 8'h07;
        13'h1C0: rddata <= 8'h3D;
        13'h1C1: rddata <= 8'h32;
        13'h1C2: rddata <= 8'h03;
        13'h1C3: rddata <= 8'hC0;
        13'h1C4: rddata <= 8'hC3;
        13'h1C5: rddata <= 8'h45;
        13'h1C6: rddata <= 8'h0F;
        13'h1C7: rddata <= 8'hCD;
        13'h1C8: rddata <= 8'hF3;
        13'h1C9: rddata <= 8'h01;
        13'h1CA: rddata <= 8'hC8;
        13'h1CB: rddata <= 8'h3E;
        13'h1CC: rddata <= 8'h15;
        13'h1CD: rddata <= 8'h32;
        13'h1CE: rddata <= 8'h03;
        13'h1CF: rddata <= 8'hC0;
        13'h1D0: rddata <= 8'hC3;
        13'h1D1: rddata <= 8'h45;
        13'h1D2: rddata <= 8'h0F;
        13'h1D3: rddata <= 8'h3A;
        13'h1D4: rddata <= 8'h03;
        13'h1D5: rddata <= 8'hC0;
        13'h1D6: rddata <= 8'hFE;
        13'h1D7: rddata <= 8'h15;
        13'h1D8: rddata <= 8'h30;
        13'h1D9: rddata <= 8'h0E;
        13'h1DA: rddata <= 8'h3C;
        13'h1DB: rddata <= 8'h47;
        13'h1DC: rddata <= 8'h3A;
        13'h1DD: rddata <= 8'h07;
        13'h1DE: rddata <= 8'hC0;
        13'h1DF: rddata <= 8'hB8;
        13'h1E0: rddata <= 8'hD8;
        13'h1E1: rddata <= 8'h78;
        13'h1E2: rddata <= 8'h32;
        13'h1E3: rddata <= 8'h03;
        13'h1E4: rddata <= 8'hC0;
        13'h1E5: rddata <= 8'hC3;
        13'h1E6: rddata <= 8'h45;
        13'h1E7: rddata <= 8'h0F;
        13'h1E8: rddata <= 8'hCD;
        13'h1E9: rddata <= 8'h03;
        13'h1EA: rddata <= 8'h02;
        13'h1EB: rddata <= 8'hC0;
        13'h1EC: rddata <= 8'hAF;
        13'h1ED: rddata <= 8'h32;
        13'h1EE: rddata <= 8'h03;
        13'h1EF: rddata <= 8'hC0;
        13'h1F0: rddata <= 8'hC3;
        13'h1F1: rddata <= 8'h45;
        13'h1F2: rddata <= 8'h0F;
        13'h1F3: rddata <= 8'h3A;
        13'h1F4: rddata <= 8'h02;
        13'h1F5: rddata <= 8'hC0;
        13'h1F6: rddata <= 8'hB7;
        13'h1F7: rddata <= 8'hC8;
        13'h1F8: rddata <= 8'h3D;
        13'h1F9: rddata <= 8'h32;
        13'h1FA: rddata <= 8'h02;
        13'h1FB: rddata <= 8'hC0;
        13'h1FC: rddata <= 8'hCD;
        13'h1FD: rddata <= 8'h27;
        13'h1FE: rddata <= 8'h02;
        13'h1FF: rddata <= 8'h3E;
        13'h200: rddata <= 8'h01;
        13'h201: rddata <= 8'hB7;
        13'h202: rddata <= 8'hC9;
        13'h203: rddata <= 8'h3A;
        13'h204: rddata <= 8'h06;
        13'h205: rddata <= 8'hC0;
        13'h206: rddata <= 8'hB7;
        13'h207: rddata <= 8'hC0;
        13'h208: rddata <= 8'h3A;
        13'h209: rddata <= 8'h02;
        13'h20A: rddata <= 8'hC0;
        13'h20B: rddata <= 8'h3C;
        13'h20C: rddata <= 8'h32;
        13'h20D: rddata <= 8'h02;
        13'h20E: rddata <= 8'hC0;
        13'h20F: rddata <= 8'hCD;
        13'h210: rddata <= 8'h27;
        13'h211: rddata <= 8'h02;
        13'h212: rddata <= 8'hAF;
        13'h213: rddata <= 8'hC9;
        13'h214: rddata <= 8'hDB;
        13'h215: rddata <= 8'hC0;
        13'h216: rddata <= 8'hEE;
        13'h217: rddata <= 8'hFF;
        13'h218: rddata <= 8'h47;
        13'h219: rddata <= 8'h3A;
        13'h21A: rddata <= 8'h04;
        13'h21B: rddata <= 8'hC0;
        13'h21C: rddata <= 8'hEE;
        13'h21D: rddata <= 8'hFF;
        13'h21E: rddata <= 8'hA0;
        13'h21F: rddata <= 8'h32;
        13'h220: rddata <= 8'h05;
        13'h221: rddata <= 8'hC0;
        13'h222: rddata <= 8'h78;
        13'h223: rddata <= 8'h32;
        13'h224: rddata <= 8'h04;
        13'h225: rddata <= 8'hC0;
        13'h226: rddata <= 8'hC9;
        13'h227: rddata <= 8'h3E;
        13'h228: rddata <= 8'h02;
        13'h229: rddata <= 8'h32;
        13'h22A: rddata <= 8'h01;
        13'h22B: rddata <= 8'hC0;
        13'h22C: rddata <= 8'hAF;
        13'h22D: rddata <= 8'h32;
        13'h22E: rddata <= 8'h00;
        13'h22F: rddata <= 8'hC0;
        13'h230: rddata <= 8'hCD;
        13'h231: rddata <= 8'h9D;
        13'h232: rddata <= 8'h0F;
        13'h233: rddata <= 8'hCD;
        13'h234: rddata <= 8'h32;
        13'h235: rddata <= 8'h10;
        13'h236: rddata <= 8'hCD;
        13'h237: rddata <= 8'h3A;
        13'h238: rddata <= 8'h10;
        13'h239: rddata <= 8'h3A;
        13'h23A: rddata <= 8'h02;
        13'h23B: rddata <= 8'hC0;
        13'h23C: rddata <= 8'h47;
        13'h23D: rddata <= 8'h04;
        13'h23E: rddata <= 8'h05;
        13'h23F: rddata <= 8'h28;
        13'h240: rddata <= 8'h0E;
        13'h241: rddata <= 8'h0E;
        13'h242: rddata <= 8'h16;
        13'h243: rddata <= 8'hC5;
        13'h244: rddata <= 8'hCD;
        13'h245: rddata <= 8'h46;
        13'h246: rddata <= 8'h10;
        13'h247: rddata <= 8'hC1;
        13'h248: rddata <= 8'h20;
        13'h249: rddata <= 8'h31;
        13'h24A: rddata <= 8'h0D;
        13'h24B: rddata <= 8'h20;
        13'h24C: rddata <= 8'hF6;
        13'h24D: rddata <= 8'h18;
        13'h24E: rddata <= 8'hEF;
        13'h24F: rddata <= 8'hAF;
        13'h250: rddata <= 8'h32;
        13'h251: rddata <= 8'h07;
        13'h252: rddata <= 8'hC0;
        13'h253: rddata <= 8'h3A;
        13'h254: rddata <= 8'h01;
        13'h255: rddata <= 8'hC0;
        13'h256: rddata <= 8'hFE;
        13'h257: rddata <= 8'h18;
        13'h258: rddata <= 8'h30;
        13'h259: rddata <= 8'h16;
        13'h25A: rddata <= 8'hCD;
        13'h25B: rddata <= 8'h46;
        13'h25C: rddata <= 8'h10;
        13'h25D: rddata <= 8'h20;
        13'h25E: rddata <= 8'h14;
        13'h25F: rddata <= 8'h3A;
        13'h260: rddata <= 8'h07;
        13'h261: rddata <= 8'hC0;
        13'h262: rddata <= 8'h3C;
        13'h263: rddata <= 8'h32;
        13'h264: rddata <= 8'h07;
        13'h265: rddata <= 8'hC0;
        13'h266: rddata <= 8'h3E;
        13'h267: rddata <= 8'h20;
        13'h268: rddata <= 8'hCD;
        13'h269: rddata <= 8'hB6;
        13'h26A: rddata <= 8'h0F;
        13'h26B: rddata <= 8'hCD;
        13'h26C: rddata <= 8'hD3;
        13'h26D: rddata <= 8'h02;
        13'h26E: rddata <= 8'h18;
        13'h26F: rddata <= 8'hE3;
        13'h270: rddata <= 8'hCD;
        13'h271: rddata <= 8'h46;
        13'h272: rddata <= 8'h10;
        13'h273: rddata <= 8'h20;
        13'h274: rddata <= 8'h06;
        13'h275: rddata <= 8'hAF;
        13'h276: rddata <= 8'h32;
        13'h277: rddata <= 8'h06;
        13'h278: rddata <= 8'hC0;
        13'h279: rddata <= 8'h18;
        13'h27A: rddata <= 8'h07;
        13'h27B: rddata <= 8'h3E;
        13'h27C: rddata <= 8'h01;
        13'h27D: rddata <= 8'h32;
        13'h27E: rddata <= 8'h06;
        13'h27F: rddata <= 8'hC0;
        13'h280: rddata <= 8'h18;
        13'h281: rddata <= 8'h00;
        13'h282: rddata <= 8'h3A;
        13'h283: rddata <= 8'h01;
        13'h284: rddata <= 8'hC0;
        13'h285: rddata <= 8'hFE;
        13'h286: rddata <= 8'h18;
        13'h287: rddata <= 8'h30;
        13'h288: rddata <= 8'h05;
        13'h289: rddata <= 8'hCD;
        13'h28A: rddata <= 8'hC7;
        13'h28B: rddata <= 8'h02;
        13'h28C: rddata <= 8'h18;
        13'h28D: rddata <= 8'hF4;
        13'h28E: rddata <= 8'h3A;
        13'h28F: rddata <= 8'h07;
        13'h290: rddata <= 8'hC0;
        13'h291: rddata <= 8'hB7;
        13'h292: rddata <= 8'h28;
        13'h293: rddata <= 8'h04;
        13'h294: rddata <= 8'hCD;
        13'h295: rddata <= 8'h45;
        13'h296: rddata <= 8'h0F;
        13'h297: rddata <= 8'hC9;
        13'h298: rddata <= 8'h3E;
        13'h299: rddata <= 8'h04;
        13'h29A: rddata <= 8'h32;
        13'h29B: rddata <= 8'h00;
        13'h29C: rddata <= 8'hC0;
        13'h29D: rddata <= 8'h3E;
        13'h29E: rddata <= 8'h08;
        13'h29F: rddata <= 8'h32;
        13'h2A0: rddata <= 8'h01;
        13'h2A1: rddata <= 8'hC0;
        13'h2A2: rddata <= 8'hCD;
        13'h2A3: rddata <= 8'h9D;
        13'h2A4: rddata <= 8'h0F;
        13'h2A5: rddata <= 8'h21;
        13'h2A6: rddata <= 8'hAF;
        13'h2A7: rddata <= 8'h02;
        13'h2A8: rddata <= 8'hCD;
        13'h2A9: rddata <= 8'hEE;
        13'h2AA: rddata <= 8'h0F;
        13'h2AB: rddata <= 8'hCD;
        13'h2AC: rddata <= 8'h7A;
        13'h2AD: rddata <= 8'h0F;
        13'h2AE: rddata <= 8'hC9;
        13'h2AF: rddata <= 8'h4E;
        13'h2B0: rddata <= 8'h6F;
        13'h2B1: rddata <= 8'h20;
        13'h2B2: rddata <= 8'h2E;
        13'h2B3: rddata <= 8'h53;
        13'h2B4: rddata <= 8'h4D;
        13'h2B5: rddata <= 8'h53;
        13'h2B6: rddata <= 8'h20;
        13'h2B7: rddata <= 8'h52;
        13'h2B8: rddata <= 8'h4F;
        13'h2B9: rddata <= 8'h4D;
        13'h2BA: rddata <= 8'h20;
        13'h2BB: rddata <= 8'h66;
        13'h2BC: rddata <= 8'h69;
        13'h2BD: rddata <= 8'h6C;
        13'h2BE: rddata <= 8'h65;
        13'h2BF: rddata <= 8'h73;
        13'h2C0: rddata <= 8'h20;
        13'h2C1: rddata <= 8'h66;
        13'h2C2: rddata <= 8'h6F;
        13'h2C3: rddata <= 8'h75;
        13'h2C4: rddata <= 8'h6E;
        13'h2C5: rddata <= 8'h64;
        13'h2C6: rddata <= 8'h00;
        13'h2C7: rddata <= 8'h3E;
        13'h2C8: rddata <= 8'h20;
        13'h2C9: rddata <= 8'hCD;
        13'h2CA: rddata <= 8'hB6;
        13'h2CB: rddata <= 8'h0F;
        13'h2CC: rddata <= 8'h3A;
        13'h2CD: rddata <= 8'h00;
        13'h2CE: rddata <= 8'hC0;
        13'h2CF: rddata <= 8'hB7;
        13'h2D0: rddata <= 8'h20;
        13'h2D1: rddata <= 8'hF5;
        13'h2D2: rddata <= 8'hC9;
        13'h2D3: rddata <= 8'h3A;
        13'h2D4: rddata <= 8'h0D;
        13'h2D5: rddata <= 8'hC0;
        13'h2D6: rddata <= 8'hCB;
        13'h2D7: rddata <= 8'h47;
        13'h2D8: rddata <= 8'h28;
        13'h2D9: rddata <= 8'h05;
        13'h2DA: rddata <= 8'h3E;
        13'h2DB: rddata <= 8'h5B;
        13'h2DC: rddata <= 8'hCD;
        13'h2DD: rddata <= 8'hB6;
        13'h2DE: rddata <= 8'h0F;
        13'h2DF: rddata <= 8'h21;
        13'h2E0: rddata <= 8'h12;
        13'h2E1: rddata <= 8'hC0;
        13'h2E2: rddata <= 8'h3A;
        13'h2E3: rddata <= 8'h08;
        13'h2E4: rddata <= 8'hC0;
        13'h2E5: rddata <= 8'h4F;
        13'h2E6: rddata <= 8'h7E;
        13'h2E7: rddata <= 8'h23;
        13'h2E8: rddata <= 8'hCD;
        13'h2E9: rddata <= 8'hB6;
        13'h2EA: rddata <= 8'h0F;
        13'h2EB: rddata <= 8'h0D;
        13'h2EC: rddata <= 8'h28;
        13'h2ED: rddata <= 8'h07;
        13'h2EE: rddata <= 8'h3A;
        13'h2EF: rddata <= 8'h00;
        13'h2F0: rddata <= 8'hC0;
        13'h2F1: rddata <= 8'hB7;
        13'h2F2: rddata <= 8'hC8;
        13'h2F3: rddata <= 8'h18;
        13'h2F4: rddata <= 8'hF1;
        13'h2F5: rddata <= 8'h3A;
        13'h2F6: rddata <= 8'h0D;
        13'h2F7: rddata <= 8'hC0;
        13'h2F8: rddata <= 8'hCB;
        13'h2F9: rddata <= 8'h47;
        13'h2FA: rddata <= 8'h28;
        13'h2FB: rddata <= 8'h05;
        13'h2FC: rddata <= 8'h3E;
        13'h2FD: rddata <= 8'h5D;
        13'h2FE: rddata <= 8'hCD;
        13'h2FF: rddata <= 8'hB6;
        13'h300: rddata <= 8'h0F;
        13'h301: rddata <= 8'h3A;
        13'h302: rddata <= 8'h00;
        13'h303: rddata <= 8'hC0;
        13'h304: rddata <= 8'hB7;
        13'h305: rddata <= 8'hC8;
        13'h306: rddata <= 8'hC3;
        13'h307: rddata <= 8'hC7;
        13'h308: rddata <= 8'h02;
        13'h309: rddata <= 8'hDB;
        13'h30A: rddata <= 8'hBF;
        13'h30B: rddata <= 8'h0E;
        13'h30C: rddata <= 8'hBF;
        13'h30D: rddata <= 8'h06;
        13'h30E: rddata <= 8'h14;
        13'h30F: rddata <= 8'h21;
        13'h310: rddata <= 8'h41;
        13'h311: rddata <= 8'h03;
        13'h312: rddata <= 8'hED;
        13'h313: rddata <= 8'hB3;
        13'h314: rddata <= 8'hAF;
        13'h315: rddata <= 8'hD3;
        13'h316: rddata <= 8'hBF;
        13'h317: rddata <= 8'h3E;
        13'h318: rddata <= 8'hC0;
        13'h319: rddata <= 8'hD3;
        13'h31A: rddata <= 8'hBF;
        13'h31B: rddata <= 8'h0E;
        13'h31C: rddata <= 8'hBE;
        13'h31D: rddata <= 8'h06;
        13'h31E: rddata <= 8'h10;
        13'h31F: rddata <= 8'h21;
        13'h320: rddata <= 8'h55;
        13'h321: rddata <= 8'h03;
        13'h322: rddata <= 8'hED;
        13'h323: rddata <= 8'hB3;
        13'h324: rddata <= 8'h06;
        13'h325: rddata <= 8'h10;
        13'h326: rddata <= 8'h21;
        13'h327: rddata <= 8'h55;
        13'h328: rddata <= 8'h03;
        13'h329: rddata <= 8'hED;
        13'h32A: rddata <= 8'hB3;
        13'h32B: rddata <= 8'hAF;
        13'h32C: rddata <= 8'hD3;
        13'h32D: rddata <= 8'hBF;
        13'h32E: rddata <= 8'h3E;
        13'h32F: rddata <= 8'h40;
        13'h330: rddata <= 8'hD3;
        13'h331: rddata <= 8'hBF;
        13'h332: rddata <= 8'h16;
        13'h333: rddata <= 8'h5F;
        13'h334: rddata <= 8'h0E;
        13'h335: rddata <= 8'hBE;
        13'h336: rddata <= 8'h21;
        13'h337: rddata <= 8'h65;
        13'h338: rddata <= 8'h03;
        13'h339: rddata <= 8'h06;
        13'h33A: rddata <= 8'h20;
        13'h33B: rddata <= 8'hED;
        13'h33C: rddata <= 8'hB3;
        13'h33D: rddata <= 8'h15;
        13'h33E: rddata <= 8'h20;
        13'h33F: rddata <= 8'hF9;
        13'h340: rddata <= 8'hC9;
        13'h341: rddata <= 8'h06;
        13'h342: rddata <= 8'h80;
        13'h343: rddata <= 8'hC0;
        13'h344: rddata <= 8'h81;
        13'h345: rddata <= 8'hFF;
        13'h346: rddata <= 8'h82;
        13'h347: rddata <= 8'hFF;
        13'h348: rddata <= 8'h83;
        13'h349: rddata <= 8'hFF;
        13'h34A: rddata <= 8'h84;
        13'h34B: rddata <= 8'hFF;
        13'h34C: rddata <= 8'h85;
        13'h34D: rddata <= 8'h00;
        13'h34E: rddata <= 8'h86;
        13'h34F: rddata <= 8'h00;
        13'h350: rddata <= 8'h87;
        13'h351: rddata <= 8'h00;
        13'h352: rddata <= 8'h88;
        13'h353: rddata <= 8'h00;
        13'h354: rddata <= 8'h89;
        13'h355: rddata <= 8'h00;
        13'h356: rddata <= 8'h03;
        13'h357: rddata <= 8'h0C;
        13'h358: rddata <= 8'h0F;
        13'h359: rddata <= 8'h30;
        13'h35A: rddata <= 8'h33;
        13'h35B: rddata <= 8'h3C;
        13'h35C: rddata <= 8'h3F;
        13'h35D: rddata <= 8'h2A;
        13'h35E: rddata <= 8'h28;
        13'h35F: rddata <= 8'h33;
        13'h360: rddata <= 8'h21;
        13'h361: rddata <= 8'h1F;
        13'h362: rddata <= 8'h1C;
        13'h363: rddata <= 8'h02;
        13'h364: rddata <= 8'h15;
        13'h365: rddata <= 8'h00;
        13'h366: rddata <= 8'h00;
        13'h367: rddata <= 8'h00;
        13'h368: rddata <= 8'h00;
        13'h369: rddata <= 8'h00;
        13'h36A: rddata <= 8'h00;
        13'h36B: rddata <= 8'h00;
        13'h36C: rddata <= 8'h00;
        13'h36D: rddata <= 8'h00;
        13'h36E: rddata <= 8'h00;
        13'h36F: rddata <= 8'h00;
        13'h370: rddata <= 8'h00;
        13'h371: rddata <= 8'h00;
        13'h372: rddata <= 8'h00;
        13'h373: rddata <= 8'h00;
        13'h374: rddata <= 8'h00;
        13'h375: rddata <= 8'h00;
        13'h376: rddata <= 8'h00;
        13'h377: rddata <= 8'h00;
        13'h378: rddata <= 8'h00;
        13'h379: rddata <= 8'h00;
        13'h37A: rddata <= 8'h00;
        13'h37B: rddata <= 8'h00;
        13'h37C: rddata <= 8'h00;
        13'h37D: rddata <= 8'h00;
        13'h37E: rddata <= 8'h00;
        13'h37F: rddata <= 8'h00;
        13'h380: rddata <= 8'h00;
        13'h381: rddata <= 8'h00;
        13'h382: rddata <= 8'h00;
        13'h383: rddata <= 8'h00;
        13'h384: rddata <= 8'h00;
        13'h385: rddata <= 8'h18;
        13'h386: rddata <= 8'h18;
        13'h387: rddata <= 8'h18;
        13'h388: rddata <= 8'h00;
        13'h389: rddata <= 8'h18;
        13'h38A: rddata <= 8'h18;
        13'h38B: rddata <= 8'h18;
        13'h38C: rddata <= 8'h00;
        13'h38D: rddata <= 8'h18;
        13'h38E: rddata <= 8'h18;
        13'h38F: rddata <= 8'h18;
        13'h390: rddata <= 8'h00;
        13'h391: rddata <= 8'h18;
        13'h392: rddata <= 8'h18;
        13'h393: rddata <= 8'h18;
        13'h394: rddata <= 8'h00;
        13'h395: rddata <= 8'h18;
        13'h396: rddata <= 8'h18;
        13'h397: rddata <= 8'h18;
        13'h398: rddata <= 8'h00;
        13'h399: rddata <= 8'h00;
        13'h39A: rddata <= 8'h00;
        13'h39B: rddata <= 8'h00;
        13'h39C: rddata <= 8'h00;
        13'h39D: rddata <= 8'h18;
        13'h39E: rddata <= 8'h18;
        13'h39F: rddata <= 8'h18;
        13'h3A0: rddata <= 8'h00;
        13'h3A1: rddata <= 8'h00;
        13'h3A2: rddata <= 8'h00;
        13'h3A3: rddata <= 8'h00;
        13'h3A4: rddata <= 8'h00;
        13'h3A5: rddata <= 8'h36;
        13'h3A6: rddata <= 8'h36;
        13'h3A7: rddata <= 8'h36;
        13'h3A8: rddata <= 8'h00;
        13'h3A9: rddata <= 8'h36;
        13'h3AA: rddata <= 8'h36;
        13'h3AB: rddata <= 8'h36;
        13'h3AC: rddata <= 8'h00;
        13'h3AD: rddata <= 8'h24;
        13'h3AE: rddata <= 8'h24;
        13'h3AF: rddata <= 8'h24;
        13'h3B0: rddata <= 8'h00;
        13'h3B1: rddata <= 8'h00;
        13'h3B2: rddata <= 8'h00;
        13'h3B3: rddata <= 8'h00;
        13'h3B4: rddata <= 8'h00;
        13'h3B5: rddata <= 8'h00;
        13'h3B6: rddata <= 8'h00;
        13'h3B7: rddata <= 8'h00;
        13'h3B8: rddata <= 8'h00;
        13'h3B9: rddata <= 8'h00;
        13'h3BA: rddata <= 8'h00;
        13'h3BB: rddata <= 8'h00;
        13'h3BC: rddata <= 8'h00;
        13'h3BD: rddata <= 8'h00;
        13'h3BE: rddata <= 8'h00;
        13'h3BF: rddata <= 8'h00;
        13'h3C0: rddata <= 8'h00;
        13'h3C1: rddata <= 8'h00;
        13'h3C2: rddata <= 8'h00;
        13'h3C3: rddata <= 8'h00;
        13'h3C4: rddata <= 8'h00;
        13'h3C5: rddata <= 8'h36;
        13'h3C6: rddata <= 8'h36;
        13'h3C7: rddata <= 8'h36;
        13'h3C8: rddata <= 8'h00;
        13'h3C9: rddata <= 8'h36;
        13'h3CA: rddata <= 8'h36;
        13'h3CB: rddata <= 8'h36;
        13'h3CC: rddata <= 8'h00;
        13'h3CD: rddata <= 8'h7F;
        13'h3CE: rddata <= 8'h7F;
        13'h3CF: rddata <= 8'h7F;
        13'h3D0: rddata <= 8'h00;
        13'h3D1: rddata <= 8'h36;
        13'h3D2: rddata <= 8'h36;
        13'h3D3: rddata <= 8'h36;
        13'h3D4: rddata <= 8'h00;
        13'h3D5: rddata <= 8'h7F;
        13'h3D6: rddata <= 8'h7F;
        13'h3D7: rddata <= 8'h7F;
        13'h3D8: rddata <= 8'h00;
        13'h3D9: rddata <= 8'h36;
        13'h3DA: rddata <= 8'h36;
        13'h3DB: rddata <= 8'h36;
        13'h3DC: rddata <= 8'h00;
        13'h3DD: rddata <= 8'h36;
        13'h3DE: rddata <= 8'h36;
        13'h3DF: rddata <= 8'h36;
        13'h3E0: rddata <= 8'h00;
        13'h3E1: rddata <= 8'h00;
        13'h3E2: rddata <= 8'h00;
        13'h3E3: rddata <= 8'h00;
        13'h3E4: rddata <= 8'h00;
        13'h3E5: rddata <= 8'h08;
        13'h3E6: rddata <= 8'h08;
        13'h3E7: rddata <= 8'h08;
        13'h3E8: rddata <= 8'h00;
        13'h3E9: rddata <= 8'h3E;
        13'h3EA: rddata <= 8'h3E;
        13'h3EB: rddata <= 8'h3E;
        13'h3EC: rddata <= 8'h00;
        13'h3ED: rddata <= 8'h68;
        13'h3EE: rddata <= 8'h68;
        13'h3EF: rddata <= 8'h68;
        13'h3F0: rddata <= 8'h00;
        13'h3F1: rddata <= 8'h3E;
        13'h3F2: rddata <= 8'h3E;
        13'h3F3: rddata <= 8'h3E;
        13'h3F4: rddata <= 8'h00;
        13'h3F5: rddata <= 8'h0B;
        13'h3F6: rddata <= 8'h0B;
        13'h3F7: rddata <= 8'h0B;
        13'h3F8: rddata <= 8'h00;
        13'h3F9: rddata <= 8'h3E;
        13'h3FA: rddata <= 8'h3E;
        13'h3FB: rddata <= 8'h3E;
        13'h3FC: rddata <= 8'h00;
        13'h3FD: rddata <= 8'h08;
        13'h3FE: rddata <= 8'h08;
        13'h3FF: rddata <= 8'h08;
        13'h400: rddata <= 8'h00;
        13'h401: rddata <= 8'h00;
        13'h402: rddata <= 8'h00;
        13'h403: rddata <= 8'h00;
        13'h404: rddata <= 8'h00;
        13'h405: rddata <= 8'h00;
        13'h406: rddata <= 8'h00;
        13'h407: rddata <= 8'h00;
        13'h408: rddata <= 8'h00;
        13'h409: rddata <= 8'h66;
        13'h40A: rddata <= 8'h66;
        13'h40B: rddata <= 8'h66;
        13'h40C: rddata <= 8'h00;
        13'h40D: rddata <= 8'h6C;
        13'h40E: rddata <= 8'h6C;
        13'h40F: rddata <= 8'h6C;
        13'h410: rddata <= 8'h00;
        13'h411: rddata <= 8'h18;
        13'h412: rddata <= 8'h18;
        13'h413: rddata <= 8'h18;
        13'h414: rddata <= 8'h00;
        13'h415: rddata <= 8'h30;
        13'h416: rddata <= 8'h30;
        13'h417: rddata <= 8'h30;
        13'h418: rddata <= 8'h00;
        13'h419: rddata <= 8'h66;
        13'h41A: rddata <= 8'h66;
        13'h41B: rddata <= 8'h66;
        13'h41C: rddata <= 8'h00;
        13'h41D: rddata <= 8'h46;
        13'h41E: rddata <= 8'h46;
        13'h41F: rddata <= 8'h46;
        13'h420: rddata <= 8'h00;
        13'h421: rddata <= 8'h00;
        13'h422: rddata <= 8'h00;
        13'h423: rddata <= 8'h00;
        13'h424: rddata <= 8'h00;
        13'h425: rddata <= 8'h1C;
        13'h426: rddata <= 8'h1C;
        13'h427: rddata <= 8'h1C;
        13'h428: rddata <= 8'h00;
        13'h429: rddata <= 8'h36;
        13'h42A: rddata <= 8'h36;
        13'h42B: rddata <= 8'h36;
        13'h42C: rddata <= 8'h00;
        13'h42D: rddata <= 8'h1C;
        13'h42E: rddata <= 8'h1C;
        13'h42F: rddata <= 8'h1C;
        13'h430: rddata <= 8'h00;
        13'h431: rddata <= 8'h3B;
        13'h432: rddata <= 8'h3B;
        13'h433: rddata <= 8'h3B;
        13'h434: rddata <= 8'h00;
        13'h435: rddata <= 8'h6E;
        13'h436: rddata <= 8'h6E;
        13'h437: rddata <= 8'h6E;
        13'h438: rddata <= 8'h00;
        13'h439: rddata <= 8'h66;
        13'h43A: rddata <= 8'h66;
        13'h43B: rddata <= 8'h66;
        13'h43C: rddata <= 8'h00;
        13'h43D: rddata <= 8'h3B;
        13'h43E: rddata <= 8'h3B;
        13'h43F: rddata <= 8'h3B;
        13'h440: rddata <= 8'h00;
        13'h441: rddata <= 8'h00;
        13'h442: rddata <= 8'h00;
        13'h443: rddata <= 8'h00;
        13'h444: rddata <= 8'h00;
        13'h445: rddata <= 8'h18;
        13'h446: rddata <= 8'h18;
        13'h447: rddata <= 8'h18;
        13'h448: rddata <= 8'h00;
        13'h449: rddata <= 8'h18;
        13'h44A: rddata <= 8'h18;
        13'h44B: rddata <= 8'h18;
        13'h44C: rddata <= 8'h00;
        13'h44D: rddata <= 8'h30;
        13'h44E: rddata <= 8'h30;
        13'h44F: rddata <= 8'h30;
        13'h450: rddata <= 8'h00;
        13'h451: rddata <= 8'h00;
        13'h452: rddata <= 8'h00;
        13'h453: rddata <= 8'h00;
        13'h454: rddata <= 8'h00;
        13'h455: rddata <= 8'h00;
        13'h456: rddata <= 8'h00;
        13'h457: rddata <= 8'h00;
        13'h458: rddata <= 8'h00;
        13'h459: rddata <= 8'h00;
        13'h45A: rddata <= 8'h00;
        13'h45B: rddata <= 8'h00;
        13'h45C: rddata <= 8'h00;
        13'h45D: rddata <= 8'h00;
        13'h45E: rddata <= 8'h00;
        13'h45F: rddata <= 8'h00;
        13'h460: rddata <= 8'h00;
        13'h461: rddata <= 8'h00;
        13'h462: rddata <= 8'h00;
        13'h463: rddata <= 8'h00;
        13'h464: rddata <= 8'h00;
        13'h465: rddata <= 8'h0C;
        13'h466: rddata <= 8'h0C;
        13'h467: rddata <= 8'h0C;
        13'h468: rddata <= 8'h00;
        13'h469: rddata <= 8'h18;
        13'h46A: rddata <= 8'h18;
        13'h46B: rddata <= 8'h18;
        13'h46C: rddata <= 8'h00;
        13'h46D: rddata <= 8'h30;
        13'h46E: rddata <= 8'h30;
        13'h46F: rddata <= 8'h30;
        13'h470: rddata <= 8'h00;
        13'h471: rddata <= 8'h30;
        13'h472: rddata <= 8'h30;
        13'h473: rddata <= 8'h30;
        13'h474: rddata <= 8'h00;
        13'h475: rddata <= 8'h30;
        13'h476: rddata <= 8'h30;
        13'h477: rddata <= 8'h30;
        13'h478: rddata <= 8'h00;
        13'h479: rddata <= 8'h18;
        13'h47A: rddata <= 8'h18;
        13'h47B: rddata <= 8'h18;
        13'h47C: rddata <= 8'h00;
        13'h47D: rddata <= 8'h0C;
        13'h47E: rddata <= 8'h0C;
        13'h47F: rddata <= 8'h0C;
        13'h480: rddata <= 8'h00;
        13'h481: rddata <= 8'h00;
        13'h482: rddata <= 8'h00;
        13'h483: rddata <= 8'h00;
        13'h484: rddata <= 8'h00;
        13'h485: rddata <= 8'h30;
        13'h486: rddata <= 8'h30;
        13'h487: rddata <= 8'h30;
        13'h488: rddata <= 8'h00;
        13'h489: rddata <= 8'h18;
        13'h48A: rddata <= 8'h18;
        13'h48B: rddata <= 8'h18;
        13'h48C: rddata <= 8'h00;
        13'h48D: rddata <= 8'h0C;
        13'h48E: rddata <= 8'h0C;
        13'h48F: rddata <= 8'h0C;
        13'h490: rddata <= 8'h00;
        13'h491: rddata <= 8'h0C;
        13'h492: rddata <= 8'h0C;
        13'h493: rddata <= 8'h0C;
        13'h494: rddata <= 8'h00;
        13'h495: rddata <= 8'h0C;
        13'h496: rddata <= 8'h0C;
        13'h497: rddata <= 8'h0C;
        13'h498: rddata <= 8'h00;
        13'h499: rddata <= 8'h18;
        13'h49A: rddata <= 8'h18;
        13'h49B: rddata <= 8'h18;
        13'h49C: rddata <= 8'h00;
        13'h49D: rddata <= 8'h30;
        13'h49E: rddata <= 8'h30;
        13'h49F: rddata <= 8'h30;
        13'h4A0: rddata <= 8'h00;
        13'h4A1: rddata <= 8'h00;
        13'h4A2: rddata <= 8'h00;
        13'h4A3: rddata <= 8'h00;
        13'h4A4: rddata <= 8'h00;
        13'h4A5: rddata <= 8'h00;
        13'h4A6: rddata <= 8'h00;
        13'h4A7: rddata <= 8'h00;
        13'h4A8: rddata <= 8'h00;
        13'h4A9: rddata <= 8'h66;
        13'h4AA: rddata <= 8'h66;
        13'h4AB: rddata <= 8'h66;
        13'h4AC: rddata <= 8'h00;
        13'h4AD: rddata <= 8'h3C;
        13'h4AE: rddata <= 8'h3C;
        13'h4AF: rddata <= 8'h3C;
        13'h4B0: rddata <= 8'h00;
        13'h4B1: rddata <= 8'hFF;
        13'h4B2: rddata <= 8'hFF;
        13'h4B3: rddata <= 8'hFF;
        13'h4B4: rddata <= 8'h00;
        13'h4B5: rddata <= 8'h3C;
        13'h4B6: rddata <= 8'h3C;
        13'h4B7: rddata <= 8'h3C;
        13'h4B8: rddata <= 8'h00;
        13'h4B9: rddata <= 8'h66;
        13'h4BA: rddata <= 8'h66;
        13'h4BB: rddata <= 8'h66;
        13'h4BC: rddata <= 8'h00;
        13'h4BD: rddata <= 8'h00;
        13'h4BE: rddata <= 8'h00;
        13'h4BF: rddata <= 8'h00;
        13'h4C0: rddata <= 8'h00;
        13'h4C1: rddata <= 8'h00;
        13'h4C2: rddata <= 8'h00;
        13'h4C3: rddata <= 8'h00;
        13'h4C4: rddata <= 8'h00;
        13'h4C5: rddata <= 8'h00;
        13'h4C6: rddata <= 8'h00;
        13'h4C7: rddata <= 8'h00;
        13'h4C8: rddata <= 8'h00;
        13'h4C9: rddata <= 8'h18;
        13'h4CA: rddata <= 8'h18;
        13'h4CB: rddata <= 8'h18;
        13'h4CC: rddata <= 8'h00;
        13'h4CD: rddata <= 8'h18;
        13'h4CE: rddata <= 8'h18;
        13'h4CF: rddata <= 8'h18;
        13'h4D0: rddata <= 8'h00;
        13'h4D1: rddata <= 8'h7E;
        13'h4D2: rddata <= 8'h7E;
        13'h4D3: rddata <= 8'h7E;
        13'h4D4: rddata <= 8'h00;
        13'h4D5: rddata <= 8'h18;
        13'h4D6: rddata <= 8'h18;
        13'h4D7: rddata <= 8'h18;
        13'h4D8: rddata <= 8'h00;
        13'h4D9: rddata <= 8'h18;
        13'h4DA: rddata <= 8'h18;
        13'h4DB: rddata <= 8'h18;
        13'h4DC: rddata <= 8'h00;
        13'h4DD: rddata <= 8'h00;
        13'h4DE: rddata <= 8'h00;
        13'h4DF: rddata <= 8'h00;
        13'h4E0: rddata <= 8'h00;
        13'h4E1: rddata <= 8'h00;
        13'h4E2: rddata <= 8'h00;
        13'h4E3: rddata <= 8'h00;
        13'h4E4: rddata <= 8'h00;
        13'h4E5: rddata <= 8'h00;
        13'h4E6: rddata <= 8'h00;
        13'h4E7: rddata <= 8'h00;
        13'h4E8: rddata <= 8'h00;
        13'h4E9: rddata <= 8'h00;
        13'h4EA: rddata <= 8'h00;
        13'h4EB: rddata <= 8'h00;
        13'h4EC: rddata <= 8'h00;
        13'h4ED: rddata <= 8'h00;
        13'h4EE: rddata <= 8'h00;
        13'h4EF: rddata <= 8'h00;
        13'h4F0: rddata <= 8'h00;
        13'h4F1: rddata <= 8'h00;
        13'h4F2: rddata <= 8'h00;
        13'h4F3: rddata <= 8'h00;
        13'h4F4: rddata <= 8'h00;
        13'h4F5: rddata <= 8'h00;
        13'h4F6: rddata <= 8'h00;
        13'h4F7: rddata <= 8'h00;
        13'h4F8: rddata <= 8'h00;
        13'h4F9: rddata <= 8'h18;
        13'h4FA: rddata <= 8'h18;
        13'h4FB: rddata <= 8'h18;
        13'h4FC: rddata <= 8'h00;
        13'h4FD: rddata <= 8'h18;
        13'h4FE: rddata <= 8'h18;
        13'h4FF: rddata <= 8'h18;
        13'h500: rddata <= 8'h00;
        13'h501: rddata <= 8'h30;
        13'h502: rddata <= 8'h30;
        13'h503: rddata <= 8'h30;
        13'h504: rddata <= 8'h00;
        13'h505: rddata <= 8'h00;
        13'h506: rddata <= 8'h00;
        13'h507: rddata <= 8'h00;
        13'h508: rddata <= 8'h00;
        13'h509: rddata <= 8'h00;
        13'h50A: rddata <= 8'h00;
        13'h50B: rddata <= 8'h00;
        13'h50C: rddata <= 8'h00;
        13'h50D: rddata <= 8'h00;
        13'h50E: rddata <= 8'h00;
        13'h50F: rddata <= 8'h00;
        13'h510: rddata <= 8'h00;
        13'h511: rddata <= 8'h3C;
        13'h512: rddata <= 8'h3C;
        13'h513: rddata <= 8'h3C;
        13'h514: rddata <= 8'h00;
        13'h515: rddata <= 8'h00;
        13'h516: rddata <= 8'h00;
        13'h517: rddata <= 8'h00;
        13'h518: rddata <= 8'h00;
        13'h519: rddata <= 8'h00;
        13'h51A: rddata <= 8'h00;
        13'h51B: rddata <= 8'h00;
        13'h51C: rddata <= 8'h00;
        13'h51D: rddata <= 8'h00;
        13'h51E: rddata <= 8'h00;
        13'h51F: rddata <= 8'h00;
        13'h520: rddata <= 8'h00;
        13'h521: rddata <= 8'h00;
        13'h522: rddata <= 8'h00;
        13'h523: rddata <= 8'h00;
        13'h524: rddata <= 8'h00;
        13'h525: rddata <= 8'h00;
        13'h526: rddata <= 8'h00;
        13'h527: rddata <= 8'h00;
        13'h528: rddata <= 8'h00;
        13'h529: rddata <= 8'h00;
        13'h52A: rddata <= 8'h00;
        13'h52B: rddata <= 8'h00;
        13'h52C: rddata <= 8'h00;
        13'h52D: rddata <= 8'h00;
        13'h52E: rddata <= 8'h00;
        13'h52F: rddata <= 8'h00;
        13'h530: rddata <= 8'h00;
        13'h531: rddata <= 8'h00;
        13'h532: rddata <= 8'h00;
        13'h533: rddata <= 8'h00;
        13'h534: rddata <= 8'h00;
        13'h535: rddata <= 8'h00;
        13'h536: rddata <= 8'h00;
        13'h537: rddata <= 8'h00;
        13'h538: rddata <= 8'h00;
        13'h539: rddata <= 8'h00;
        13'h53A: rddata <= 8'h00;
        13'h53B: rddata <= 8'h00;
        13'h53C: rddata <= 8'h00;
        13'h53D: rddata <= 8'h18;
        13'h53E: rddata <= 8'h18;
        13'h53F: rddata <= 8'h18;
        13'h540: rddata <= 8'h00;
        13'h541: rddata <= 8'h00;
        13'h542: rddata <= 8'h00;
        13'h543: rddata <= 8'h00;
        13'h544: rddata <= 8'h00;
        13'h545: rddata <= 8'h02;
        13'h546: rddata <= 8'h02;
        13'h547: rddata <= 8'h02;
        13'h548: rddata <= 8'h00;
        13'h549: rddata <= 8'h06;
        13'h54A: rddata <= 8'h06;
        13'h54B: rddata <= 8'h06;
        13'h54C: rddata <= 8'h00;
        13'h54D: rddata <= 8'h0C;
        13'h54E: rddata <= 8'h0C;
        13'h54F: rddata <= 8'h0C;
        13'h550: rddata <= 8'h00;
        13'h551: rddata <= 8'h18;
        13'h552: rddata <= 8'h18;
        13'h553: rddata <= 8'h18;
        13'h554: rddata <= 8'h00;
        13'h555: rddata <= 8'h30;
        13'h556: rddata <= 8'h30;
        13'h557: rddata <= 8'h30;
        13'h558: rddata <= 8'h00;
        13'h559: rddata <= 8'h60;
        13'h55A: rddata <= 8'h60;
        13'h55B: rddata <= 8'h60;
        13'h55C: rddata <= 8'h00;
        13'h55D: rddata <= 8'h40;
        13'h55E: rddata <= 8'h40;
        13'h55F: rddata <= 8'h40;
        13'h560: rddata <= 8'h00;
        13'h561: rddata <= 8'h00;
        13'h562: rddata <= 8'h00;
        13'h563: rddata <= 8'h00;
        13'h564: rddata <= 8'h00;
        13'h565: rddata <= 8'h1C;
        13'h566: rddata <= 8'h1C;
        13'h567: rddata <= 8'h1C;
        13'h568: rddata <= 8'h00;
        13'h569: rddata <= 8'h26;
        13'h56A: rddata <= 8'h26;
        13'h56B: rddata <= 8'h26;
        13'h56C: rddata <= 8'h00;
        13'h56D: rddata <= 8'h63;
        13'h56E: rddata <= 8'h63;
        13'h56F: rddata <= 8'h63;
        13'h570: rddata <= 8'h00;
        13'h571: rddata <= 8'h63;
        13'h572: rddata <= 8'h63;
        13'h573: rddata <= 8'h63;
        13'h574: rddata <= 8'h00;
        13'h575: rddata <= 8'h63;
        13'h576: rddata <= 8'h63;
        13'h577: rddata <= 8'h63;
        13'h578: rddata <= 8'h00;
        13'h579: rddata <= 8'h32;
        13'h57A: rddata <= 8'h32;
        13'h57B: rddata <= 8'h32;
        13'h57C: rddata <= 8'h00;
        13'h57D: rddata <= 8'h1C;
        13'h57E: rddata <= 8'h1C;
        13'h57F: rddata <= 8'h1C;
        13'h580: rddata <= 8'h00;
        13'h581: rddata <= 8'h00;
        13'h582: rddata <= 8'h00;
        13'h583: rddata <= 8'h00;
        13'h584: rddata <= 8'h00;
        13'h585: rddata <= 8'h0C;
        13'h586: rddata <= 8'h0C;
        13'h587: rddata <= 8'h0C;
        13'h588: rddata <= 8'h00;
        13'h589: rddata <= 8'h1C;
        13'h58A: rddata <= 8'h1C;
        13'h58B: rddata <= 8'h1C;
        13'h58C: rddata <= 8'h00;
        13'h58D: rddata <= 8'h0C;
        13'h58E: rddata <= 8'h0C;
        13'h58F: rddata <= 8'h0C;
        13'h590: rddata <= 8'h00;
        13'h591: rddata <= 8'h0C;
        13'h592: rddata <= 8'h0C;
        13'h593: rddata <= 8'h0C;
        13'h594: rddata <= 8'h00;
        13'h595: rddata <= 8'h0C;
        13'h596: rddata <= 8'h0C;
        13'h597: rddata <= 8'h0C;
        13'h598: rddata <= 8'h00;
        13'h599: rddata <= 8'h0C;
        13'h59A: rddata <= 8'h0C;
        13'h59B: rddata <= 8'h0C;
        13'h59C: rddata <= 8'h00;
        13'h59D: rddata <= 8'h3F;
        13'h59E: rddata <= 8'h3F;
        13'h59F: rddata <= 8'h3F;
        13'h5A0: rddata <= 8'h00;
        13'h5A1: rddata <= 8'h00;
        13'h5A2: rddata <= 8'h00;
        13'h5A3: rddata <= 8'h00;
        13'h5A4: rddata <= 8'h00;
        13'h5A5: rddata <= 8'h3E;
        13'h5A6: rddata <= 8'h3E;
        13'h5A7: rddata <= 8'h3E;
        13'h5A8: rddata <= 8'h00;
        13'h5A9: rddata <= 8'h63;
        13'h5AA: rddata <= 8'h63;
        13'h5AB: rddata <= 8'h63;
        13'h5AC: rddata <= 8'h00;
        13'h5AD: rddata <= 8'h07;
        13'h5AE: rddata <= 8'h07;
        13'h5AF: rddata <= 8'h07;
        13'h5B0: rddata <= 8'h00;
        13'h5B1: rddata <= 8'h1E;
        13'h5B2: rddata <= 8'h1E;
        13'h5B3: rddata <= 8'h1E;
        13'h5B4: rddata <= 8'h00;
        13'h5B5: rddata <= 8'h3C;
        13'h5B6: rddata <= 8'h3C;
        13'h5B7: rddata <= 8'h3C;
        13'h5B8: rddata <= 8'h00;
        13'h5B9: rddata <= 8'h70;
        13'h5BA: rddata <= 8'h70;
        13'h5BB: rddata <= 8'h70;
        13'h5BC: rddata <= 8'h00;
        13'h5BD: rddata <= 8'h7F;
        13'h5BE: rddata <= 8'h7F;
        13'h5BF: rddata <= 8'h7F;
        13'h5C0: rddata <= 8'h00;
        13'h5C1: rddata <= 8'h00;
        13'h5C2: rddata <= 8'h00;
        13'h5C3: rddata <= 8'h00;
        13'h5C4: rddata <= 8'h00;
        13'h5C5: rddata <= 8'h3F;
        13'h5C6: rddata <= 8'h3F;
        13'h5C7: rddata <= 8'h3F;
        13'h5C8: rddata <= 8'h00;
        13'h5C9: rddata <= 8'h06;
        13'h5CA: rddata <= 8'h06;
        13'h5CB: rddata <= 8'h06;
        13'h5CC: rddata <= 8'h00;
        13'h5CD: rddata <= 8'h0C;
        13'h5CE: rddata <= 8'h0C;
        13'h5CF: rddata <= 8'h0C;
        13'h5D0: rddata <= 8'h00;
        13'h5D1: rddata <= 8'h1E;
        13'h5D2: rddata <= 8'h1E;
        13'h5D3: rddata <= 8'h1E;
        13'h5D4: rddata <= 8'h00;
        13'h5D5: rddata <= 8'h03;
        13'h5D6: rddata <= 8'h03;
        13'h5D7: rddata <= 8'h03;
        13'h5D8: rddata <= 8'h00;
        13'h5D9: rddata <= 8'h63;
        13'h5DA: rddata <= 8'h63;
        13'h5DB: rddata <= 8'h63;
        13'h5DC: rddata <= 8'h00;
        13'h5DD: rddata <= 8'h3E;
        13'h5DE: rddata <= 8'h3E;
        13'h5DF: rddata <= 8'h3E;
        13'h5E0: rddata <= 8'h00;
        13'h5E1: rddata <= 8'h00;
        13'h5E2: rddata <= 8'h00;
        13'h5E3: rddata <= 8'h00;
        13'h5E4: rddata <= 8'h00;
        13'h5E5: rddata <= 8'h06;
        13'h5E6: rddata <= 8'h06;
        13'h5E7: rddata <= 8'h06;
        13'h5E8: rddata <= 8'h00;
        13'h5E9: rddata <= 8'h0E;
        13'h5EA: rddata <= 8'h0E;
        13'h5EB: rddata <= 8'h0E;
        13'h5EC: rddata <= 8'h00;
        13'h5ED: rddata <= 8'h1E;
        13'h5EE: rddata <= 8'h1E;
        13'h5EF: rddata <= 8'h1E;
        13'h5F0: rddata <= 8'h00;
        13'h5F1: rddata <= 8'h36;
        13'h5F2: rddata <= 8'h36;
        13'h5F3: rddata <= 8'h36;
        13'h5F4: rddata <= 8'h00;
        13'h5F5: rddata <= 8'h66;
        13'h5F6: rddata <= 8'h66;
        13'h5F7: rddata <= 8'h66;
        13'h5F8: rddata <= 8'h00;
        13'h5F9: rddata <= 8'h7F;
        13'h5FA: rddata <= 8'h7F;
        13'h5FB: rddata <= 8'h7F;
        13'h5FC: rddata <= 8'h00;
        13'h5FD: rddata <= 8'h06;
        13'h5FE: rddata <= 8'h06;
        13'h5FF: rddata <= 8'h06;
        13'h600: rddata <= 8'h00;
        13'h601: rddata <= 8'h00;
        13'h602: rddata <= 8'h00;
        13'h603: rddata <= 8'h00;
        13'h604: rddata <= 8'h00;
        13'h605: rddata <= 8'h7E;
        13'h606: rddata <= 8'h7E;
        13'h607: rddata <= 8'h7E;
        13'h608: rddata <= 8'h00;
        13'h609: rddata <= 8'h60;
        13'h60A: rddata <= 8'h60;
        13'h60B: rddata <= 8'h60;
        13'h60C: rddata <= 8'h00;
        13'h60D: rddata <= 8'h7E;
        13'h60E: rddata <= 8'h7E;
        13'h60F: rddata <= 8'h7E;
        13'h610: rddata <= 8'h00;
        13'h611: rddata <= 8'h03;
        13'h612: rddata <= 8'h03;
        13'h613: rddata <= 8'h03;
        13'h614: rddata <= 8'h00;
        13'h615: rddata <= 8'h03;
        13'h616: rddata <= 8'h03;
        13'h617: rddata <= 8'h03;
        13'h618: rddata <= 8'h00;
        13'h619: rddata <= 8'h63;
        13'h61A: rddata <= 8'h63;
        13'h61B: rddata <= 8'h63;
        13'h61C: rddata <= 8'h00;
        13'h61D: rddata <= 8'h3E;
        13'h61E: rddata <= 8'h3E;
        13'h61F: rddata <= 8'h3E;
        13'h620: rddata <= 8'h00;
        13'h621: rddata <= 8'h00;
        13'h622: rddata <= 8'h00;
        13'h623: rddata <= 8'h00;
        13'h624: rddata <= 8'h00;
        13'h625: rddata <= 8'h1E;
        13'h626: rddata <= 8'h1E;
        13'h627: rddata <= 8'h1E;
        13'h628: rddata <= 8'h00;
        13'h629: rddata <= 8'h30;
        13'h62A: rddata <= 8'h30;
        13'h62B: rddata <= 8'h30;
        13'h62C: rddata <= 8'h00;
        13'h62D: rddata <= 8'h60;
        13'h62E: rddata <= 8'h60;
        13'h62F: rddata <= 8'h60;
        13'h630: rddata <= 8'h00;
        13'h631: rddata <= 8'h7E;
        13'h632: rddata <= 8'h7E;
        13'h633: rddata <= 8'h7E;
        13'h634: rddata <= 8'h00;
        13'h635: rddata <= 8'h63;
        13'h636: rddata <= 8'h63;
        13'h637: rddata <= 8'h63;
        13'h638: rddata <= 8'h00;
        13'h639: rddata <= 8'h63;
        13'h63A: rddata <= 8'h63;
        13'h63B: rddata <= 8'h63;
        13'h63C: rddata <= 8'h00;
        13'h63D: rddata <= 8'h3E;
        13'h63E: rddata <= 8'h3E;
        13'h63F: rddata <= 8'h3E;
        13'h640: rddata <= 8'h00;
        13'h641: rddata <= 8'h00;
        13'h642: rddata <= 8'h00;
        13'h643: rddata <= 8'h00;
        13'h644: rddata <= 8'h00;
        13'h645: rddata <= 8'h7F;
        13'h646: rddata <= 8'h7F;
        13'h647: rddata <= 8'h7F;
        13'h648: rddata <= 8'h00;
        13'h649: rddata <= 8'h63;
        13'h64A: rddata <= 8'h63;
        13'h64B: rddata <= 8'h63;
        13'h64C: rddata <= 8'h00;
        13'h64D: rddata <= 8'h06;
        13'h64E: rddata <= 8'h06;
        13'h64F: rddata <= 8'h06;
        13'h650: rddata <= 8'h00;
        13'h651: rddata <= 8'h0C;
        13'h652: rddata <= 8'h0C;
        13'h653: rddata <= 8'h0C;
        13'h654: rddata <= 8'h00;
        13'h655: rddata <= 8'h18;
        13'h656: rddata <= 8'h18;
        13'h657: rddata <= 8'h18;
        13'h658: rddata <= 8'h00;
        13'h659: rddata <= 8'h18;
        13'h65A: rddata <= 8'h18;
        13'h65B: rddata <= 8'h18;
        13'h65C: rddata <= 8'h00;
        13'h65D: rddata <= 8'h18;
        13'h65E: rddata <= 8'h18;
        13'h65F: rddata <= 8'h18;
        13'h660: rddata <= 8'h00;
        13'h661: rddata <= 8'h00;
        13'h662: rddata <= 8'h00;
        13'h663: rddata <= 8'h00;
        13'h664: rddata <= 8'h00;
        13'h665: rddata <= 8'h3C;
        13'h666: rddata <= 8'h3C;
        13'h667: rddata <= 8'h3C;
        13'h668: rddata <= 8'h00;
        13'h669: rddata <= 8'h62;
        13'h66A: rddata <= 8'h62;
        13'h66B: rddata <= 8'h62;
        13'h66C: rddata <= 8'h00;
        13'h66D: rddata <= 8'h72;
        13'h66E: rddata <= 8'h72;
        13'h66F: rddata <= 8'h72;
        13'h670: rddata <= 8'h00;
        13'h671: rddata <= 8'h3C;
        13'h672: rddata <= 8'h3C;
        13'h673: rddata <= 8'h3C;
        13'h674: rddata <= 8'h00;
        13'h675: rddata <= 8'h4F;
        13'h676: rddata <= 8'h4F;
        13'h677: rddata <= 8'h4F;
        13'h678: rddata <= 8'h00;
        13'h679: rddata <= 8'h43;
        13'h67A: rddata <= 8'h43;
        13'h67B: rddata <= 8'h43;
        13'h67C: rddata <= 8'h00;
        13'h67D: rddata <= 8'h3E;
        13'h67E: rddata <= 8'h3E;
        13'h67F: rddata <= 8'h3E;
        13'h680: rddata <= 8'h00;
        13'h681: rddata <= 8'h00;
        13'h682: rddata <= 8'h00;
        13'h683: rddata <= 8'h00;
        13'h684: rddata <= 8'h00;
        13'h685: rddata <= 8'h3E;
        13'h686: rddata <= 8'h3E;
        13'h687: rddata <= 8'h3E;
        13'h688: rddata <= 8'h00;
        13'h689: rddata <= 8'h63;
        13'h68A: rddata <= 8'h63;
        13'h68B: rddata <= 8'h63;
        13'h68C: rddata <= 8'h00;
        13'h68D: rddata <= 8'h63;
        13'h68E: rddata <= 8'h63;
        13'h68F: rddata <= 8'h63;
        13'h690: rddata <= 8'h00;
        13'h691: rddata <= 8'h3F;
        13'h692: rddata <= 8'h3F;
        13'h693: rddata <= 8'h3F;
        13'h694: rddata <= 8'h00;
        13'h695: rddata <= 8'h03;
        13'h696: rddata <= 8'h03;
        13'h697: rddata <= 8'h03;
        13'h698: rddata <= 8'h00;
        13'h699: rddata <= 8'h06;
        13'h69A: rddata <= 8'h06;
        13'h69B: rddata <= 8'h06;
        13'h69C: rddata <= 8'h00;
        13'h69D: rddata <= 8'h3C;
        13'h69E: rddata <= 8'h3C;
        13'h69F: rddata <= 8'h3C;
        13'h6A0: rddata <= 8'h00;
        13'h6A1: rddata <= 8'h00;
        13'h6A2: rddata <= 8'h00;
        13'h6A3: rddata <= 8'h00;
        13'h6A4: rddata <= 8'h00;
        13'h6A5: rddata <= 8'h00;
        13'h6A6: rddata <= 8'h00;
        13'h6A7: rddata <= 8'h00;
        13'h6A8: rddata <= 8'h00;
        13'h6A9: rddata <= 8'h00;
        13'h6AA: rddata <= 8'h00;
        13'h6AB: rddata <= 8'h00;
        13'h6AC: rddata <= 8'h00;
        13'h6AD: rddata <= 8'h00;
        13'h6AE: rddata <= 8'h00;
        13'h6AF: rddata <= 8'h00;
        13'h6B0: rddata <= 8'h00;
        13'h6B1: rddata <= 8'h18;
        13'h6B2: rddata <= 8'h18;
        13'h6B3: rddata <= 8'h18;
        13'h6B4: rddata <= 8'h00;
        13'h6B5: rddata <= 8'h00;
        13'h6B6: rddata <= 8'h00;
        13'h6B7: rddata <= 8'h00;
        13'h6B8: rddata <= 8'h00;
        13'h6B9: rddata <= 8'h18;
        13'h6BA: rddata <= 8'h18;
        13'h6BB: rddata <= 8'h18;
        13'h6BC: rddata <= 8'h00;
        13'h6BD: rddata <= 8'h00;
        13'h6BE: rddata <= 8'h00;
        13'h6BF: rddata <= 8'h00;
        13'h6C0: rddata <= 8'h00;
        13'h6C1: rddata <= 8'h00;
        13'h6C2: rddata <= 8'h00;
        13'h6C3: rddata <= 8'h00;
        13'h6C4: rddata <= 8'h00;
        13'h6C5: rddata <= 8'h00;
        13'h6C6: rddata <= 8'h00;
        13'h6C7: rddata <= 8'h00;
        13'h6C8: rddata <= 8'h00;
        13'h6C9: rddata <= 8'h00;
        13'h6CA: rddata <= 8'h00;
        13'h6CB: rddata <= 8'h00;
        13'h6CC: rddata <= 8'h00;
        13'h6CD: rddata <= 8'h00;
        13'h6CE: rddata <= 8'h00;
        13'h6CF: rddata <= 8'h00;
        13'h6D0: rddata <= 8'h00;
        13'h6D1: rddata <= 8'h18;
        13'h6D2: rddata <= 8'h18;
        13'h6D3: rddata <= 8'h18;
        13'h6D4: rddata <= 8'h00;
        13'h6D5: rddata <= 8'h00;
        13'h6D6: rddata <= 8'h00;
        13'h6D7: rddata <= 8'h00;
        13'h6D8: rddata <= 8'h00;
        13'h6D9: rddata <= 8'h18;
        13'h6DA: rddata <= 8'h18;
        13'h6DB: rddata <= 8'h18;
        13'h6DC: rddata <= 8'h00;
        13'h6DD: rddata <= 8'h18;
        13'h6DE: rddata <= 8'h18;
        13'h6DF: rddata <= 8'h18;
        13'h6E0: rddata <= 8'h00;
        13'h6E1: rddata <= 8'h30;
        13'h6E2: rddata <= 8'h30;
        13'h6E3: rddata <= 8'h30;
        13'h6E4: rddata <= 8'h00;
        13'h6E5: rddata <= 8'h00;
        13'h6E6: rddata <= 8'h00;
        13'h6E7: rddata <= 8'h00;
        13'h6E8: rddata <= 8'h00;
        13'h6E9: rddata <= 8'h00;
        13'h6EA: rddata <= 8'h00;
        13'h6EB: rddata <= 8'h00;
        13'h6EC: rddata <= 8'h00;
        13'h6ED: rddata <= 8'h0C;
        13'h6EE: rddata <= 8'h0C;
        13'h6EF: rddata <= 8'h0C;
        13'h6F0: rddata <= 8'h00;
        13'h6F1: rddata <= 8'h18;
        13'h6F2: rddata <= 8'h18;
        13'h6F3: rddata <= 8'h18;
        13'h6F4: rddata <= 8'h00;
        13'h6F5: rddata <= 8'h30;
        13'h6F6: rddata <= 8'h30;
        13'h6F7: rddata <= 8'h30;
        13'h6F8: rddata <= 8'h00;
        13'h6F9: rddata <= 8'h18;
        13'h6FA: rddata <= 8'h18;
        13'h6FB: rddata <= 8'h18;
        13'h6FC: rddata <= 8'h00;
        13'h6FD: rddata <= 8'h0C;
        13'h6FE: rddata <= 8'h0C;
        13'h6FF: rddata <= 8'h0C;
        13'h700: rddata <= 8'h00;
        13'h701: rddata <= 8'h00;
        13'h702: rddata <= 8'h00;
        13'h703: rddata <= 8'h00;
        13'h704: rddata <= 8'h00;
        13'h705: rddata <= 8'h00;
        13'h706: rddata <= 8'h00;
        13'h707: rddata <= 8'h00;
        13'h708: rddata <= 8'h00;
        13'h709: rddata <= 8'h00;
        13'h70A: rddata <= 8'h00;
        13'h70B: rddata <= 8'h00;
        13'h70C: rddata <= 8'h00;
        13'h70D: rddata <= 8'h00;
        13'h70E: rddata <= 8'h00;
        13'h70F: rddata <= 8'h00;
        13'h710: rddata <= 8'h00;
        13'h711: rddata <= 8'h3E;
        13'h712: rddata <= 8'h3E;
        13'h713: rddata <= 8'h3E;
        13'h714: rddata <= 8'h00;
        13'h715: rddata <= 8'h00;
        13'h716: rddata <= 8'h00;
        13'h717: rddata <= 8'h00;
        13'h718: rddata <= 8'h00;
        13'h719: rddata <= 8'h3E;
        13'h71A: rddata <= 8'h3E;
        13'h71B: rddata <= 8'h3E;
        13'h71C: rddata <= 8'h00;
        13'h71D: rddata <= 8'h00;
        13'h71E: rddata <= 8'h00;
        13'h71F: rddata <= 8'h00;
        13'h720: rddata <= 8'h00;
        13'h721: rddata <= 8'h00;
        13'h722: rddata <= 8'h00;
        13'h723: rddata <= 8'h00;
        13'h724: rddata <= 8'h00;
        13'h725: rddata <= 8'h00;
        13'h726: rddata <= 8'h00;
        13'h727: rddata <= 8'h00;
        13'h728: rddata <= 8'h00;
        13'h729: rddata <= 8'h00;
        13'h72A: rddata <= 8'h00;
        13'h72B: rddata <= 8'h00;
        13'h72C: rddata <= 8'h00;
        13'h72D: rddata <= 8'h30;
        13'h72E: rddata <= 8'h30;
        13'h72F: rddata <= 8'h30;
        13'h730: rddata <= 8'h00;
        13'h731: rddata <= 8'h18;
        13'h732: rddata <= 8'h18;
        13'h733: rddata <= 8'h18;
        13'h734: rddata <= 8'h00;
        13'h735: rddata <= 8'h0C;
        13'h736: rddata <= 8'h0C;
        13'h737: rddata <= 8'h0C;
        13'h738: rddata <= 8'h00;
        13'h739: rddata <= 8'h18;
        13'h73A: rddata <= 8'h18;
        13'h73B: rddata <= 8'h18;
        13'h73C: rddata <= 8'h00;
        13'h73D: rddata <= 8'h30;
        13'h73E: rddata <= 8'h30;
        13'h73F: rddata <= 8'h30;
        13'h740: rddata <= 8'h00;
        13'h741: rddata <= 8'h00;
        13'h742: rddata <= 8'h00;
        13'h743: rddata <= 8'h00;
        13'h744: rddata <= 8'h00;
        13'h745: rddata <= 8'h3C;
        13'h746: rddata <= 8'h3C;
        13'h747: rddata <= 8'h3C;
        13'h748: rddata <= 8'h00;
        13'h749: rddata <= 8'h66;
        13'h74A: rddata <= 8'h66;
        13'h74B: rddata <= 8'h66;
        13'h74C: rddata <= 8'h00;
        13'h74D: rddata <= 8'h06;
        13'h74E: rddata <= 8'h06;
        13'h74F: rddata <= 8'h06;
        13'h750: rddata <= 8'h00;
        13'h751: rddata <= 8'h0C;
        13'h752: rddata <= 8'h0C;
        13'h753: rddata <= 8'h0C;
        13'h754: rddata <= 8'h00;
        13'h755: rddata <= 8'h18;
        13'h756: rddata <= 8'h18;
        13'h757: rddata <= 8'h18;
        13'h758: rddata <= 8'h00;
        13'h759: rddata <= 8'h00;
        13'h75A: rddata <= 8'h00;
        13'h75B: rddata <= 8'h00;
        13'h75C: rddata <= 8'h00;
        13'h75D: rddata <= 8'h18;
        13'h75E: rddata <= 8'h18;
        13'h75F: rddata <= 8'h18;
        13'h760: rddata <= 8'h00;
        13'h761: rddata <= 8'h00;
        13'h762: rddata <= 8'h00;
        13'h763: rddata <= 8'h00;
        13'h764: rddata <= 8'h00;
        13'h765: rddata <= 8'h3E;
        13'h766: rddata <= 8'h3E;
        13'h767: rddata <= 8'h3E;
        13'h768: rddata <= 8'h00;
        13'h769: rddata <= 8'h63;
        13'h76A: rddata <= 8'h63;
        13'h76B: rddata <= 8'h63;
        13'h76C: rddata <= 8'h00;
        13'h76D: rddata <= 8'h6F;
        13'h76E: rddata <= 8'h6F;
        13'h76F: rddata <= 8'h6F;
        13'h770: rddata <= 8'h00;
        13'h771: rddata <= 8'h6B;
        13'h772: rddata <= 8'h6B;
        13'h773: rddata <= 8'h6B;
        13'h774: rddata <= 8'h00;
        13'h775: rddata <= 8'h6E;
        13'h776: rddata <= 8'h6E;
        13'h777: rddata <= 8'h6E;
        13'h778: rddata <= 8'h00;
        13'h779: rddata <= 8'h60;
        13'h77A: rddata <= 8'h60;
        13'h77B: rddata <= 8'h60;
        13'h77C: rddata <= 8'h00;
        13'h77D: rddata <= 8'h3E;
        13'h77E: rddata <= 8'h3E;
        13'h77F: rddata <= 8'h3E;
        13'h780: rddata <= 8'h00;
        13'h781: rddata <= 8'h00;
        13'h782: rddata <= 8'h00;
        13'h783: rddata <= 8'h00;
        13'h784: rddata <= 8'h00;
        13'h785: rddata <= 8'h18;
        13'h786: rddata <= 8'h18;
        13'h787: rddata <= 8'h18;
        13'h788: rddata <= 8'h00;
        13'h789: rddata <= 8'h3C;
        13'h78A: rddata <= 8'h3C;
        13'h78B: rddata <= 8'h3C;
        13'h78C: rddata <= 8'h00;
        13'h78D: rddata <= 8'h66;
        13'h78E: rddata <= 8'h66;
        13'h78F: rddata <= 8'h66;
        13'h790: rddata <= 8'h00;
        13'h791: rddata <= 8'h66;
        13'h792: rddata <= 8'h66;
        13'h793: rddata <= 8'h66;
        13'h794: rddata <= 8'h00;
        13'h795: rddata <= 8'h7E;
        13'h796: rddata <= 8'h7E;
        13'h797: rddata <= 8'h7E;
        13'h798: rddata <= 8'h00;
        13'h799: rddata <= 8'h66;
        13'h79A: rddata <= 8'h66;
        13'h79B: rddata <= 8'h66;
        13'h79C: rddata <= 8'h00;
        13'h79D: rddata <= 8'h66;
        13'h79E: rddata <= 8'h66;
        13'h79F: rddata <= 8'h66;
        13'h7A0: rddata <= 8'h00;
        13'h7A1: rddata <= 8'h00;
        13'h7A2: rddata <= 8'h00;
        13'h7A3: rddata <= 8'h00;
        13'h7A4: rddata <= 8'h00;
        13'h7A5: rddata <= 8'h7C;
        13'h7A6: rddata <= 8'h7C;
        13'h7A7: rddata <= 8'h7C;
        13'h7A8: rddata <= 8'h00;
        13'h7A9: rddata <= 8'h66;
        13'h7AA: rddata <= 8'h66;
        13'h7AB: rddata <= 8'h66;
        13'h7AC: rddata <= 8'h00;
        13'h7AD: rddata <= 8'h66;
        13'h7AE: rddata <= 8'h66;
        13'h7AF: rddata <= 8'h66;
        13'h7B0: rddata <= 8'h00;
        13'h7B1: rddata <= 8'h7C;
        13'h7B2: rddata <= 8'h7C;
        13'h7B3: rddata <= 8'h7C;
        13'h7B4: rddata <= 8'h00;
        13'h7B5: rddata <= 8'h66;
        13'h7B6: rddata <= 8'h66;
        13'h7B7: rddata <= 8'h66;
        13'h7B8: rddata <= 8'h00;
        13'h7B9: rddata <= 8'h66;
        13'h7BA: rddata <= 8'h66;
        13'h7BB: rddata <= 8'h66;
        13'h7BC: rddata <= 8'h00;
        13'h7BD: rddata <= 8'h7C;
        13'h7BE: rddata <= 8'h7C;
        13'h7BF: rddata <= 8'h7C;
        13'h7C0: rddata <= 8'h00;
        13'h7C1: rddata <= 8'h00;
        13'h7C2: rddata <= 8'h00;
        13'h7C3: rddata <= 8'h00;
        13'h7C4: rddata <= 8'h00;
        13'h7C5: rddata <= 8'h3C;
        13'h7C6: rddata <= 8'h3C;
        13'h7C7: rddata <= 8'h3C;
        13'h7C8: rddata <= 8'h00;
        13'h7C9: rddata <= 8'h66;
        13'h7CA: rddata <= 8'h66;
        13'h7CB: rddata <= 8'h66;
        13'h7CC: rddata <= 8'h00;
        13'h7CD: rddata <= 8'h60;
        13'h7CE: rddata <= 8'h60;
        13'h7CF: rddata <= 8'h60;
        13'h7D0: rddata <= 8'h00;
        13'h7D1: rddata <= 8'h60;
        13'h7D2: rddata <= 8'h60;
        13'h7D3: rddata <= 8'h60;
        13'h7D4: rddata <= 8'h00;
        13'h7D5: rddata <= 8'h60;
        13'h7D6: rddata <= 8'h60;
        13'h7D7: rddata <= 8'h60;
        13'h7D8: rddata <= 8'h00;
        13'h7D9: rddata <= 8'h66;
        13'h7DA: rddata <= 8'h66;
        13'h7DB: rddata <= 8'h66;
        13'h7DC: rddata <= 8'h00;
        13'h7DD: rddata <= 8'h3C;
        13'h7DE: rddata <= 8'h3C;
        13'h7DF: rddata <= 8'h3C;
        13'h7E0: rddata <= 8'h00;
        13'h7E1: rddata <= 8'h00;
        13'h7E2: rddata <= 8'h00;
        13'h7E3: rddata <= 8'h00;
        13'h7E4: rddata <= 8'h00;
        13'h7E5: rddata <= 8'h7C;
        13'h7E6: rddata <= 8'h7C;
        13'h7E7: rddata <= 8'h7C;
        13'h7E8: rddata <= 8'h00;
        13'h7E9: rddata <= 8'h66;
        13'h7EA: rddata <= 8'h66;
        13'h7EB: rddata <= 8'h66;
        13'h7EC: rddata <= 8'h00;
        13'h7ED: rddata <= 8'h66;
        13'h7EE: rddata <= 8'h66;
        13'h7EF: rddata <= 8'h66;
        13'h7F0: rddata <= 8'h00;
        13'h7F1: rddata <= 8'h66;
        13'h7F2: rddata <= 8'h66;
        13'h7F3: rddata <= 8'h66;
        13'h7F4: rddata <= 8'h00;
        13'h7F5: rddata <= 8'h66;
        13'h7F6: rddata <= 8'h66;
        13'h7F7: rddata <= 8'h66;
        13'h7F8: rddata <= 8'h00;
        13'h7F9: rddata <= 8'h66;
        13'h7FA: rddata <= 8'h66;
        13'h7FB: rddata <= 8'h66;
        13'h7FC: rddata <= 8'h00;
        13'h7FD: rddata <= 8'h7C;
        13'h7FE: rddata <= 8'h7C;
        13'h7FF: rddata <= 8'h7C;
        13'h800: rddata <= 8'h00;
        13'h801: rddata <= 8'h00;
        13'h802: rddata <= 8'h00;
        13'h803: rddata <= 8'h00;
        13'h804: rddata <= 8'h00;
        13'h805: rddata <= 8'h7E;
        13'h806: rddata <= 8'h7E;
        13'h807: rddata <= 8'h7E;
        13'h808: rddata <= 8'h00;
        13'h809: rddata <= 8'h60;
        13'h80A: rddata <= 8'h60;
        13'h80B: rddata <= 8'h60;
        13'h80C: rddata <= 8'h00;
        13'h80D: rddata <= 8'h60;
        13'h80E: rddata <= 8'h60;
        13'h80F: rddata <= 8'h60;
        13'h810: rddata <= 8'h00;
        13'h811: rddata <= 8'h78;
        13'h812: rddata <= 8'h78;
        13'h813: rddata <= 8'h78;
        13'h814: rddata <= 8'h00;
        13'h815: rddata <= 8'h60;
        13'h816: rddata <= 8'h60;
        13'h817: rddata <= 8'h60;
        13'h818: rddata <= 8'h00;
        13'h819: rddata <= 8'h60;
        13'h81A: rddata <= 8'h60;
        13'h81B: rddata <= 8'h60;
        13'h81C: rddata <= 8'h00;
        13'h81D: rddata <= 8'h7E;
        13'h81E: rddata <= 8'h7E;
        13'h81F: rddata <= 8'h7E;
        13'h820: rddata <= 8'h00;
        13'h821: rddata <= 8'h00;
        13'h822: rddata <= 8'h00;
        13'h823: rddata <= 8'h00;
        13'h824: rddata <= 8'h00;
        13'h825: rddata <= 8'h7E;
        13'h826: rddata <= 8'h7E;
        13'h827: rddata <= 8'h7E;
        13'h828: rddata <= 8'h00;
        13'h829: rddata <= 8'h60;
        13'h82A: rddata <= 8'h60;
        13'h82B: rddata <= 8'h60;
        13'h82C: rddata <= 8'h00;
        13'h82D: rddata <= 8'h60;
        13'h82E: rddata <= 8'h60;
        13'h82F: rddata <= 8'h60;
        13'h830: rddata <= 8'h00;
        13'h831: rddata <= 8'h78;
        13'h832: rddata <= 8'h78;
        13'h833: rddata <= 8'h78;
        13'h834: rddata <= 8'h00;
        13'h835: rddata <= 8'h60;
        13'h836: rddata <= 8'h60;
        13'h837: rddata <= 8'h60;
        13'h838: rddata <= 8'h00;
        13'h839: rddata <= 8'h60;
        13'h83A: rddata <= 8'h60;
        13'h83B: rddata <= 8'h60;
        13'h83C: rddata <= 8'h00;
        13'h83D: rddata <= 8'h60;
        13'h83E: rddata <= 8'h60;
        13'h83F: rddata <= 8'h60;
        13'h840: rddata <= 8'h00;
        13'h841: rddata <= 8'h00;
        13'h842: rddata <= 8'h00;
        13'h843: rddata <= 8'h00;
        13'h844: rddata <= 8'h00;
        13'h845: rddata <= 8'h3C;
        13'h846: rddata <= 8'h3C;
        13'h847: rddata <= 8'h3C;
        13'h848: rddata <= 8'h00;
        13'h849: rddata <= 8'h66;
        13'h84A: rddata <= 8'h66;
        13'h84B: rddata <= 8'h66;
        13'h84C: rddata <= 8'h00;
        13'h84D: rddata <= 8'h60;
        13'h84E: rddata <= 8'h60;
        13'h84F: rddata <= 8'h60;
        13'h850: rddata <= 8'h00;
        13'h851: rddata <= 8'h6E;
        13'h852: rddata <= 8'h6E;
        13'h853: rddata <= 8'h6E;
        13'h854: rddata <= 8'h00;
        13'h855: rddata <= 8'h66;
        13'h856: rddata <= 8'h66;
        13'h857: rddata <= 8'h66;
        13'h858: rddata <= 8'h00;
        13'h859: rddata <= 8'h66;
        13'h85A: rddata <= 8'h66;
        13'h85B: rddata <= 8'h66;
        13'h85C: rddata <= 8'h00;
        13'h85D: rddata <= 8'h3C;
        13'h85E: rddata <= 8'h3C;
        13'h85F: rddata <= 8'h3C;
        13'h860: rddata <= 8'h00;
        13'h861: rddata <= 8'h00;
        13'h862: rddata <= 8'h00;
        13'h863: rddata <= 8'h00;
        13'h864: rddata <= 8'h00;
        13'h865: rddata <= 8'h66;
        13'h866: rddata <= 8'h66;
        13'h867: rddata <= 8'h66;
        13'h868: rddata <= 8'h00;
        13'h869: rddata <= 8'h66;
        13'h86A: rddata <= 8'h66;
        13'h86B: rddata <= 8'h66;
        13'h86C: rddata <= 8'h00;
        13'h86D: rddata <= 8'h66;
        13'h86E: rddata <= 8'h66;
        13'h86F: rddata <= 8'h66;
        13'h870: rddata <= 8'h00;
        13'h871: rddata <= 8'h7E;
        13'h872: rddata <= 8'h7E;
        13'h873: rddata <= 8'h7E;
        13'h874: rddata <= 8'h00;
        13'h875: rddata <= 8'h66;
        13'h876: rddata <= 8'h66;
        13'h877: rddata <= 8'h66;
        13'h878: rddata <= 8'h00;
        13'h879: rddata <= 8'h66;
        13'h87A: rddata <= 8'h66;
        13'h87B: rddata <= 8'h66;
        13'h87C: rddata <= 8'h00;
        13'h87D: rddata <= 8'h66;
        13'h87E: rddata <= 8'h66;
        13'h87F: rddata <= 8'h66;
        13'h880: rddata <= 8'h00;
        13'h881: rddata <= 8'h00;
        13'h882: rddata <= 8'h00;
        13'h883: rddata <= 8'h00;
        13'h884: rddata <= 8'h00;
        13'h885: rddata <= 8'h3C;
        13'h886: rddata <= 8'h3C;
        13'h887: rddata <= 8'h3C;
        13'h888: rddata <= 8'h00;
        13'h889: rddata <= 8'h18;
        13'h88A: rddata <= 8'h18;
        13'h88B: rddata <= 8'h18;
        13'h88C: rddata <= 8'h00;
        13'h88D: rddata <= 8'h18;
        13'h88E: rddata <= 8'h18;
        13'h88F: rddata <= 8'h18;
        13'h890: rddata <= 8'h00;
        13'h891: rddata <= 8'h18;
        13'h892: rddata <= 8'h18;
        13'h893: rddata <= 8'h18;
        13'h894: rddata <= 8'h00;
        13'h895: rddata <= 8'h18;
        13'h896: rddata <= 8'h18;
        13'h897: rddata <= 8'h18;
        13'h898: rddata <= 8'h00;
        13'h899: rddata <= 8'h18;
        13'h89A: rddata <= 8'h18;
        13'h89B: rddata <= 8'h18;
        13'h89C: rddata <= 8'h00;
        13'h89D: rddata <= 8'h3C;
        13'h89E: rddata <= 8'h3C;
        13'h89F: rddata <= 8'h3C;
        13'h8A0: rddata <= 8'h00;
        13'h8A1: rddata <= 8'h00;
        13'h8A2: rddata <= 8'h00;
        13'h8A3: rddata <= 8'h00;
        13'h8A4: rddata <= 8'h00;
        13'h8A5: rddata <= 8'h00;
        13'h8A6: rddata <= 8'h00;
        13'h8A7: rddata <= 8'h00;
        13'h8A8: rddata <= 8'h00;
        13'h8A9: rddata <= 8'h06;
        13'h8AA: rddata <= 8'h06;
        13'h8AB: rddata <= 8'h06;
        13'h8AC: rddata <= 8'h00;
        13'h8AD: rddata <= 8'h06;
        13'h8AE: rddata <= 8'h06;
        13'h8AF: rddata <= 8'h06;
        13'h8B0: rddata <= 8'h00;
        13'h8B1: rddata <= 8'h06;
        13'h8B2: rddata <= 8'h06;
        13'h8B3: rddata <= 8'h06;
        13'h8B4: rddata <= 8'h00;
        13'h8B5: rddata <= 8'h06;
        13'h8B6: rddata <= 8'h06;
        13'h8B7: rddata <= 8'h06;
        13'h8B8: rddata <= 8'h00;
        13'h8B9: rddata <= 8'h66;
        13'h8BA: rddata <= 8'h66;
        13'h8BB: rddata <= 8'h66;
        13'h8BC: rddata <= 8'h00;
        13'h8BD: rddata <= 8'h3C;
        13'h8BE: rddata <= 8'h3C;
        13'h8BF: rddata <= 8'h3C;
        13'h8C0: rddata <= 8'h00;
        13'h8C1: rddata <= 8'h00;
        13'h8C2: rddata <= 8'h00;
        13'h8C3: rddata <= 8'h00;
        13'h8C4: rddata <= 8'h00;
        13'h8C5: rddata <= 8'h02;
        13'h8C6: rddata <= 8'h02;
        13'h8C7: rddata <= 8'h02;
        13'h8C8: rddata <= 8'h00;
        13'h8C9: rddata <= 8'h66;
        13'h8CA: rddata <= 8'h66;
        13'h8CB: rddata <= 8'h66;
        13'h8CC: rddata <= 8'h00;
        13'h8CD: rddata <= 8'h6C;
        13'h8CE: rddata <= 8'h6C;
        13'h8CF: rddata <= 8'h6C;
        13'h8D0: rddata <= 8'h00;
        13'h8D1: rddata <= 8'h78;
        13'h8D2: rddata <= 8'h78;
        13'h8D3: rddata <= 8'h78;
        13'h8D4: rddata <= 8'h00;
        13'h8D5: rddata <= 8'h6C;
        13'h8D6: rddata <= 8'h6C;
        13'h8D7: rddata <= 8'h6C;
        13'h8D8: rddata <= 8'h00;
        13'h8D9: rddata <= 8'h66;
        13'h8DA: rddata <= 8'h66;
        13'h8DB: rddata <= 8'h66;
        13'h8DC: rddata <= 8'h00;
        13'h8DD: rddata <= 8'h66;
        13'h8DE: rddata <= 8'h66;
        13'h8DF: rddata <= 8'h66;
        13'h8E0: rddata <= 8'h00;
        13'h8E1: rddata <= 8'h00;
        13'h8E2: rddata <= 8'h00;
        13'h8E3: rddata <= 8'h00;
        13'h8E4: rddata <= 8'h00;
        13'h8E5: rddata <= 8'h60;
        13'h8E6: rddata <= 8'h60;
        13'h8E7: rddata <= 8'h60;
        13'h8E8: rddata <= 8'h00;
        13'h8E9: rddata <= 8'h60;
        13'h8EA: rddata <= 8'h60;
        13'h8EB: rddata <= 8'h60;
        13'h8EC: rddata <= 8'h00;
        13'h8ED: rddata <= 8'h60;
        13'h8EE: rddata <= 8'h60;
        13'h8EF: rddata <= 8'h60;
        13'h8F0: rddata <= 8'h00;
        13'h8F1: rddata <= 8'h60;
        13'h8F2: rddata <= 8'h60;
        13'h8F3: rddata <= 8'h60;
        13'h8F4: rddata <= 8'h00;
        13'h8F5: rddata <= 8'h60;
        13'h8F6: rddata <= 8'h60;
        13'h8F7: rddata <= 8'h60;
        13'h8F8: rddata <= 8'h00;
        13'h8F9: rddata <= 8'h60;
        13'h8FA: rddata <= 8'h60;
        13'h8FB: rddata <= 8'h60;
        13'h8FC: rddata <= 8'h00;
        13'h8FD: rddata <= 8'h7E;
        13'h8FE: rddata <= 8'h7E;
        13'h8FF: rddata <= 8'h7E;
        13'h900: rddata <= 8'h00;
        13'h901: rddata <= 8'h00;
        13'h902: rddata <= 8'h00;
        13'h903: rddata <= 8'h00;
        13'h904: rddata <= 8'h00;
        13'h905: rddata <= 8'hC6;
        13'h906: rddata <= 8'hC6;
        13'h907: rddata <= 8'hC6;
        13'h908: rddata <= 8'h00;
        13'h909: rddata <= 8'hEE;
        13'h90A: rddata <= 8'hEE;
        13'h90B: rddata <= 8'hEE;
        13'h90C: rddata <= 8'h00;
        13'h90D: rddata <= 8'hFE;
        13'h90E: rddata <= 8'hFE;
        13'h90F: rddata <= 8'hFE;
        13'h910: rddata <= 8'h00;
        13'h911: rddata <= 8'hD6;
        13'h912: rddata <= 8'hD6;
        13'h913: rddata <= 8'hD6;
        13'h914: rddata <= 8'h00;
        13'h915: rddata <= 8'hC6;
        13'h916: rddata <= 8'hC6;
        13'h917: rddata <= 8'hC6;
        13'h918: rddata <= 8'h00;
        13'h919: rddata <= 8'hC6;
        13'h91A: rddata <= 8'hC6;
        13'h91B: rddata <= 8'hC6;
        13'h91C: rddata <= 8'h00;
        13'h91D: rddata <= 8'hC6;
        13'h91E: rddata <= 8'hC6;
        13'h91F: rddata <= 8'hC6;
        13'h920: rddata <= 8'h00;
        13'h921: rddata <= 8'h00;
        13'h922: rddata <= 8'h00;
        13'h923: rddata <= 8'h00;
        13'h924: rddata <= 8'h00;
        13'h925: rddata <= 8'h66;
        13'h926: rddata <= 8'h66;
        13'h927: rddata <= 8'h66;
        13'h928: rddata <= 8'h00;
        13'h929: rddata <= 8'h76;
        13'h92A: rddata <= 8'h76;
        13'h92B: rddata <= 8'h76;
        13'h92C: rddata <= 8'h00;
        13'h92D: rddata <= 8'h7E;
        13'h92E: rddata <= 8'h7E;
        13'h92F: rddata <= 8'h7E;
        13'h930: rddata <= 8'h00;
        13'h931: rddata <= 8'h6E;
        13'h932: rddata <= 8'h6E;
        13'h933: rddata <= 8'h6E;
        13'h934: rddata <= 8'h00;
        13'h935: rddata <= 8'h66;
        13'h936: rddata <= 8'h66;
        13'h937: rddata <= 8'h66;
        13'h938: rddata <= 8'h00;
        13'h939: rddata <= 8'h66;
        13'h93A: rddata <= 8'h66;
        13'h93B: rddata <= 8'h66;
        13'h93C: rddata <= 8'h00;
        13'h93D: rddata <= 8'h66;
        13'h93E: rddata <= 8'h66;
        13'h93F: rddata <= 8'h66;
        13'h940: rddata <= 8'h00;
        13'h941: rddata <= 8'h00;
        13'h942: rddata <= 8'h00;
        13'h943: rddata <= 8'h00;
        13'h944: rddata <= 8'h00;
        13'h945: rddata <= 8'h3C;
        13'h946: rddata <= 8'h3C;
        13'h947: rddata <= 8'h3C;
        13'h948: rddata <= 8'h00;
        13'h949: rddata <= 8'h66;
        13'h94A: rddata <= 8'h66;
        13'h94B: rddata <= 8'h66;
        13'h94C: rddata <= 8'h00;
        13'h94D: rddata <= 8'h66;
        13'h94E: rddata <= 8'h66;
        13'h94F: rddata <= 8'h66;
        13'h950: rddata <= 8'h00;
        13'h951: rddata <= 8'h66;
        13'h952: rddata <= 8'h66;
        13'h953: rddata <= 8'h66;
        13'h954: rddata <= 8'h00;
        13'h955: rddata <= 8'h66;
        13'h956: rddata <= 8'h66;
        13'h957: rddata <= 8'h66;
        13'h958: rddata <= 8'h00;
        13'h959: rddata <= 8'h66;
        13'h95A: rddata <= 8'h66;
        13'h95B: rddata <= 8'h66;
        13'h95C: rddata <= 8'h00;
        13'h95D: rddata <= 8'h3C;
        13'h95E: rddata <= 8'h3C;
        13'h95F: rddata <= 8'h3C;
        13'h960: rddata <= 8'h00;
        13'h961: rddata <= 8'h00;
        13'h962: rddata <= 8'h00;
        13'h963: rddata <= 8'h00;
        13'h964: rddata <= 8'h00;
        13'h965: rddata <= 8'h7C;
        13'h966: rddata <= 8'h7C;
        13'h967: rddata <= 8'h7C;
        13'h968: rddata <= 8'h00;
        13'h969: rddata <= 8'h66;
        13'h96A: rddata <= 8'h66;
        13'h96B: rddata <= 8'h66;
        13'h96C: rddata <= 8'h00;
        13'h96D: rddata <= 8'h66;
        13'h96E: rddata <= 8'h66;
        13'h96F: rddata <= 8'h66;
        13'h970: rddata <= 8'h00;
        13'h971: rddata <= 8'h7C;
        13'h972: rddata <= 8'h7C;
        13'h973: rddata <= 8'h7C;
        13'h974: rddata <= 8'h00;
        13'h975: rddata <= 8'h60;
        13'h976: rddata <= 8'h60;
        13'h977: rddata <= 8'h60;
        13'h978: rddata <= 8'h00;
        13'h979: rddata <= 8'h60;
        13'h97A: rddata <= 8'h60;
        13'h97B: rddata <= 8'h60;
        13'h97C: rddata <= 8'h00;
        13'h97D: rddata <= 8'h60;
        13'h97E: rddata <= 8'h60;
        13'h97F: rddata <= 8'h60;
        13'h980: rddata <= 8'h00;
        13'h981: rddata <= 8'h00;
        13'h982: rddata <= 8'h00;
        13'h983: rddata <= 8'h00;
        13'h984: rddata <= 8'h00;
        13'h985: rddata <= 8'h3C;
        13'h986: rddata <= 8'h3C;
        13'h987: rddata <= 8'h3C;
        13'h988: rddata <= 8'h00;
        13'h989: rddata <= 8'h66;
        13'h98A: rddata <= 8'h66;
        13'h98B: rddata <= 8'h66;
        13'h98C: rddata <= 8'h00;
        13'h98D: rddata <= 8'h66;
        13'h98E: rddata <= 8'h66;
        13'h98F: rddata <= 8'h66;
        13'h990: rddata <= 8'h00;
        13'h991: rddata <= 8'h66;
        13'h992: rddata <= 8'h66;
        13'h993: rddata <= 8'h66;
        13'h994: rddata <= 8'h00;
        13'h995: rddata <= 8'h66;
        13'h996: rddata <= 8'h66;
        13'h997: rddata <= 8'h66;
        13'h998: rddata <= 8'h00;
        13'h999: rddata <= 8'h6E;
        13'h99A: rddata <= 8'h6E;
        13'h99B: rddata <= 8'h6E;
        13'h99C: rddata <= 8'h00;
        13'h99D: rddata <= 8'h3C;
        13'h99E: rddata <= 8'h3C;
        13'h99F: rddata <= 8'h3C;
        13'h9A0: rddata <= 8'h00;
        13'h9A1: rddata <= 8'h06;
        13'h9A2: rddata <= 8'h06;
        13'h9A3: rddata <= 8'h06;
        13'h9A4: rddata <= 8'h00;
        13'h9A5: rddata <= 8'h7C;
        13'h9A6: rddata <= 8'h7C;
        13'h9A7: rddata <= 8'h7C;
        13'h9A8: rddata <= 8'h00;
        13'h9A9: rddata <= 8'h66;
        13'h9AA: rddata <= 8'h66;
        13'h9AB: rddata <= 8'h66;
        13'h9AC: rddata <= 8'h00;
        13'h9AD: rddata <= 8'h66;
        13'h9AE: rddata <= 8'h66;
        13'h9AF: rddata <= 8'h66;
        13'h9B0: rddata <= 8'h00;
        13'h9B1: rddata <= 8'h7C;
        13'h9B2: rddata <= 8'h7C;
        13'h9B3: rddata <= 8'h7C;
        13'h9B4: rddata <= 8'h00;
        13'h9B5: rddata <= 8'h66;
        13'h9B6: rddata <= 8'h66;
        13'h9B7: rddata <= 8'h66;
        13'h9B8: rddata <= 8'h00;
        13'h9B9: rddata <= 8'h66;
        13'h9BA: rddata <= 8'h66;
        13'h9BB: rddata <= 8'h66;
        13'h9BC: rddata <= 8'h00;
        13'h9BD: rddata <= 8'h66;
        13'h9BE: rddata <= 8'h66;
        13'h9BF: rddata <= 8'h66;
        13'h9C0: rddata <= 8'h00;
        13'h9C1: rddata <= 8'h00;
        13'h9C2: rddata <= 8'h00;
        13'h9C3: rddata <= 8'h00;
        13'h9C4: rddata <= 8'h00;
        13'h9C5: rddata <= 8'h3C;
        13'h9C6: rddata <= 8'h3C;
        13'h9C7: rddata <= 8'h3C;
        13'h9C8: rddata <= 8'h00;
        13'h9C9: rddata <= 8'h66;
        13'h9CA: rddata <= 8'h66;
        13'h9CB: rddata <= 8'h66;
        13'h9CC: rddata <= 8'h00;
        13'h9CD: rddata <= 8'h60;
        13'h9CE: rddata <= 8'h60;
        13'h9CF: rddata <= 8'h60;
        13'h9D0: rddata <= 8'h00;
        13'h9D1: rddata <= 8'h3C;
        13'h9D2: rddata <= 8'h3C;
        13'h9D3: rddata <= 8'h3C;
        13'h9D4: rddata <= 8'h00;
        13'h9D5: rddata <= 8'h06;
        13'h9D6: rddata <= 8'h06;
        13'h9D7: rddata <= 8'h06;
        13'h9D8: rddata <= 8'h00;
        13'h9D9: rddata <= 8'h66;
        13'h9DA: rddata <= 8'h66;
        13'h9DB: rddata <= 8'h66;
        13'h9DC: rddata <= 8'h00;
        13'h9DD: rddata <= 8'h3C;
        13'h9DE: rddata <= 8'h3C;
        13'h9DF: rddata <= 8'h3C;
        13'h9E0: rddata <= 8'h00;
        13'h9E1: rddata <= 8'h00;
        13'h9E2: rddata <= 8'h00;
        13'h9E3: rddata <= 8'h00;
        13'h9E4: rddata <= 8'h00;
        13'h9E5: rddata <= 8'h7E;
        13'h9E6: rddata <= 8'h7E;
        13'h9E7: rddata <= 8'h7E;
        13'h9E8: rddata <= 8'h00;
        13'h9E9: rddata <= 8'h18;
        13'h9EA: rddata <= 8'h18;
        13'h9EB: rddata <= 8'h18;
        13'h9EC: rddata <= 8'h00;
        13'h9ED: rddata <= 8'h18;
        13'h9EE: rddata <= 8'h18;
        13'h9EF: rddata <= 8'h18;
        13'h9F0: rddata <= 8'h00;
        13'h9F1: rddata <= 8'h18;
        13'h9F2: rddata <= 8'h18;
        13'h9F3: rddata <= 8'h18;
        13'h9F4: rddata <= 8'h00;
        13'h9F5: rddata <= 8'h18;
        13'h9F6: rddata <= 8'h18;
        13'h9F7: rddata <= 8'h18;
        13'h9F8: rddata <= 8'h00;
        13'h9F9: rddata <= 8'h18;
        13'h9FA: rddata <= 8'h18;
        13'h9FB: rddata <= 8'h18;
        13'h9FC: rddata <= 8'h00;
        13'h9FD: rddata <= 8'h18;
        13'h9FE: rddata <= 8'h18;
        13'h9FF: rddata <= 8'h18;
        13'hA00: rddata <= 8'h00;
        13'hA01: rddata <= 8'h00;
        13'hA02: rddata <= 8'h00;
        13'hA03: rddata <= 8'h00;
        13'hA04: rddata <= 8'h00;
        13'hA05: rddata <= 8'h66;
        13'hA06: rddata <= 8'h66;
        13'hA07: rddata <= 8'h66;
        13'hA08: rddata <= 8'h00;
        13'hA09: rddata <= 8'h66;
        13'hA0A: rddata <= 8'h66;
        13'hA0B: rddata <= 8'h66;
        13'hA0C: rddata <= 8'h00;
        13'hA0D: rddata <= 8'h66;
        13'hA0E: rddata <= 8'h66;
        13'hA0F: rddata <= 8'h66;
        13'hA10: rddata <= 8'h00;
        13'hA11: rddata <= 8'h66;
        13'hA12: rddata <= 8'h66;
        13'hA13: rddata <= 8'h66;
        13'hA14: rddata <= 8'h00;
        13'hA15: rddata <= 8'h66;
        13'hA16: rddata <= 8'h66;
        13'hA17: rddata <= 8'h66;
        13'hA18: rddata <= 8'h00;
        13'hA19: rddata <= 8'h66;
        13'hA1A: rddata <= 8'h66;
        13'hA1B: rddata <= 8'h66;
        13'hA1C: rddata <= 8'h00;
        13'hA1D: rddata <= 8'h3C;
        13'hA1E: rddata <= 8'h3C;
        13'hA1F: rddata <= 8'h3C;
        13'hA20: rddata <= 8'h00;
        13'hA21: rddata <= 8'h00;
        13'hA22: rddata <= 8'h00;
        13'hA23: rddata <= 8'h00;
        13'hA24: rddata <= 8'h00;
        13'hA25: rddata <= 8'h66;
        13'hA26: rddata <= 8'h66;
        13'hA27: rddata <= 8'h66;
        13'hA28: rddata <= 8'h00;
        13'hA29: rddata <= 8'h66;
        13'hA2A: rddata <= 8'h66;
        13'hA2B: rddata <= 8'h66;
        13'hA2C: rddata <= 8'h00;
        13'hA2D: rddata <= 8'h66;
        13'hA2E: rddata <= 8'h66;
        13'hA2F: rddata <= 8'h66;
        13'hA30: rddata <= 8'h00;
        13'hA31: rddata <= 8'h66;
        13'hA32: rddata <= 8'h66;
        13'hA33: rddata <= 8'h66;
        13'hA34: rddata <= 8'h00;
        13'hA35: rddata <= 8'h66;
        13'hA36: rddata <= 8'h66;
        13'hA37: rddata <= 8'h66;
        13'hA38: rddata <= 8'h00;
        13'hA39: rddata <= 8'h3C;
        13'hA3A: rddata <= 8'h3C;
        13'hA3B: rddata <= 8'h3C;
        13'hA3C: rddata <= 8'h00;
        13'hA3D: rddata <= 8'h18;
        13'hA3E: rddata <= 8'h18;
        13'hA3F: rddata <= 8'h18;
        13'hA40: rddata <= 8'h00;
        13'hA41: rddata <= 8'h00;
        13'hA42: rddata <= 8'h00;
        13'hA43: rddata <= 8'h00;
        13'hA44: rddata <= 8'h00;
        13'hA45: rddata <= 8'hC6;
        13'hA46: rddata <= 8'hC6;
        13'hA47: rddata <= 8'hC6;
        13'hA48: rddata <= 8'h00;
        13'hA49: rddata <= 8'hC6;
        13'hA4A: rddata <= 8'hC6;
        13'hA4B: rddata <= 8'hC6;
        13'hA4C: rddata <= 8'h00;
        13'hA4D: rddata <= 8'hC6;
        13'hA4E: rddata <= 8'hC6;
        13'hA4F: rddata <= 8'hC6;
        13'hA50: rddata <= 8'h00;
        13'hA51: rddata <= 8'hD6;
        13'hA52: rddata <= 8'hD6;
        13'hA53: rddata <= 8'hD6;
        13'hA54: rddata <= 8'h00;
        13'hA55: rddata <= 8'hD6;
        13'hA56: rddata <= 8'hD6;
        13'hA57: rddata <= 8'hD6;
        13'hA58: rddata <= 8'h00;
        13'hA59: rddata <= 8'hFE;
        13'hA5A: rddata <= 8'hFE;
        13'hA5B: rddata <= 8'hFE;
        13'hA5C: rddata <= 8'h00;
        13'hA5D: rddata <= 8'h6C;
        13'hA5E: rddata <= 8'h6C;
        13'hA5F: rddata <= 8'h6C;
        13'hA60: rddata <= 8'h00;
        13'hA61: rddata <= 8'h00;
        13'hA62: rddata <= 8'h00;
        13'hA63: rddata <= 8'h00;
        13'hA64: rddata <= 8'h00;
        13'hA65: rddata <= 8'h66;
        13'hA66: rddata <= 8'h66;
        13'hA67: rddata <= 8'h66;
        13'hA68: rddata <= 8'h00;
        13'hA69: rddata <= 8'h66;
        13'hA6A: rddata <= 8'h66;
        13'hA6B: rddata <= 8'h66;
        13'hA6C: rddata <= 8'h00;
        13'hA6D: rddata <= 8'h3C;
        13'hA6E: rddata <= 8'h3C;
        13'hA6F: rddata <= 8'h3C;
        13'hA70: rddata <= 8'h00;
        13'hA71: rddata <= 8'h18;
        13'hA72: rddata <= 8'h18;
        13'hA73: rddata <= 8'h18;
        13'hA74: rddata <= 8'h00;
        13'hA75: rddata <= 8'h3C;
        13'hA76: rddata <= 8'h3C;
        13'hA77: rddata <= 8'h3C;
        13'hA78: rddata <= 8'h00;
        13'hA79: rddata <= 8'h66;
        13'hA7A: rddata <= 8'h66;
        13'hA7B: rddata <= 8'h66;
        13'hA7C: rddata <= 8'h00;
        13'hA7D: rddata <= 8'h66;
        13'hA7E: rddata <= 8'h66;
        13'hA7F: rddata <= 8'h66;
        13'hA80: rddata <= 8'h00;
        13'hA81: rddata <= 8'h00;
        13'hA82: rddata <= 8'h00;
        13'hA83: rddata <= 8'h00;
        13'hA84: rddata <= 8'h00;
        13'hA85: rddata <= 8'h66;
        13'hA86: rddata <= 8'h66;
        13'hA87: rddata <= 8'h66;
        13'hA88: rddata <= 8'h00;
        13'hA89: rddata <= 8'h66;
        13'hA8A: rddata <= 8'h66;
        13'hA8B: rddata <= 8'h66;
        13'hA8C: rddata <= 8'h00;
        13'hA8D: rddata <= 8'h66;
        13'hA8E: rddata <= 8'h66;
        13'hA8F: rddata <= 8'h66;
        13'hA90: rddata <= 8'h00;
        13'hA91: rddata <= 8'h3C;
        13'hA92: rddata <= 8'h3C;
        13'hA93: rddata <= 8'h3C;
        13'hA94: rddata <= 8'h00;
        13'hA95: rddata <= 8'h18;
        13'hA96: rddata <= 8'h18;
        13'hA97: rddata <= 8'h18;
        13'hA98: rddata <= 8'h00;
        13'hA99: rddata <= 8'h18;
        13'hA9A: rddata <= 8'h18;
        13'hA9B: rddata <= 8'h18;
        13'hA9C: rddata <= 8'h00;
        13'hA9D: rddata <= 8'h18;
        13'hA9E: rddata <= 8'h18;
        13'hA9F: rddata <= 8'h18;
        13'hAA0: rddata <= 8'h00;
        13'hAA1: rddata <= 8'h00;
        13'hAA2: rddata <= 8'h00;
        13'hAA3: rddata <= 8'h00;
        13'hAA4: rddata <= 8'h00;
        13'hAA5: rddata <= 8'h7E;
        13'hAA6: rddata <= 8'h7E;
        13'hAA7: rddata <= 8'h7E;
        13'hAA8: rddata <= 8'h00;
        13'hAA9: rddata <= 8'h06;
        13'hAAA: rddata <= 8'h06;
        13'hAAB: rddata <= 8'h06;
        13'hAAC: rddata <= 8'h00;
        13'hAAD: rddata <= 8'h0C;
        13'hAAE: rddata <= 8'h0C;
        13'hAAF: rddata <= 8'h0C;
        13'hAB0: rddata <= 8'h00;
        13'hAB1: rddata <= 8'h18;
        13'hAB2: rddata <= 8'h18;
        13'hAB3: rddata <= 8'h18;
        13'hAB4: rddata <= 8'h00;
        13'hAB5: rddata <= 8'h30;
        13'hAB6: rddata <= 8'h30;
        13'hAB7: rddata <= 8'h30;
        13'hAB8: rddata <= 8'h00;
        13'hAB9: rddata <= 8'h60;
        13'hABA: rddata <= 8'h60;
        13'hABB: rddata <= 8'h60;
        13'hABC: rddata <= 8'h00;
        13'hABD: rddata <= 8'h7E;
        13'hABE: rddata <= 8'h7E;
        13'hABF: rddata <= 8'h7E;
        13'hAC0: rddata <= 8'h00;
        13'hAC1: rddata <= 8'h00;
        13'hAC2: rddata <= 8'h00;
        13'hAC3: rddata <= 8'h00;
        13'hAC4: rddata <= 8'h00;
        13'hAC5: rddata <= 8'h3C;
        13'hAC6: rddata <= 8'h3C;
        13'hAC7: rddata <= 8'h3C;
        13'hAC8: rddata <= 8'h00;
        13'hAC9: rddata <= 8'h30;
        13'hACA: rddata <= 8'h30;
        13'hACB: rddata <= 8'h30;
        13'hACC: rddata <= 8'h00;
        13'hACD: rddata <= 8'h30;
        13'hACE: rddata <= 8'h30;
        13'hACF: rddata <= 8'h30;
        13'hAD0: rddata <= 8'h00;
        13'hAD1: rddata <= 8'h30;
        13'hAD2: rddata <= 8'h30;
        13'hAD3: rddata <= 8'h30;
        13'hAD4: rddata <= 8'h00;
        13'hAD5: rddata <= 8'h30;
        13'hAD6: rddata <= 8'h30;
        13'hAD7: rddata <= 8'h30;
        13'hAD8: rddata <= 8'h00;
        13'hAD9: rddata <= 8'h30;
        13'hADA: rddata <= 8'h30;
        13'hADB: rddata <= 8'h30;
        13'hADC: rddata <= 8'h00;
        13'hADD: rddata <= 8'h3C;
        13'hADE: rddata <= 8'h3C;
        13'hADF: rddata <= 8'h3C;
        13'hAE0: rddata <= 8'h00;
        13'hAE1: rddata <= 8'h00;
        13'hAE2: rddata <= 8'h00;
        13'hAE3: rddata <= 8'h00;
        13'hAE4: rddata <= 8'h00;
        13'hAE5: rddata <= 8'h40;
        13'hAE6: rddata <= 8'h40;
        13'hAE7: rddata <= 8'h40;
        13'hAE8: rddata <= 8'h00;
        13'hAE9: rddata <= 8'h60;
        13'hAEA: rddata <= 8'h60;
        13'hAEB: rddata <= 8'h60;
        13'hAEC: rddata <= 8'h00;
        13'hAED: rddata <= 8'h30;
        13'hAEE: rddata <= 8'h30;
        13'hAEF: rddata <= 8'h30;
        13'hAF0: rddata <= 8'h00;
        13'hAF1: rddata <= 8'h18;
        13'hAF2: rddata <= 8'h18;
        13'hAF3: rddata <= 8'h18;
        13'hAF4: rddata <= 8'h00;
        13'hAF5: rddata <= 8'h0C;
        13'hAF6: rddata <= 8'h0C;
        13'hAF7: rddata <= 8'h0C;
        13'hAF8: rddata <= 8'h00;
        13'hAF9: rddata <= 8'h06;
        13'hAFA: rddata <= 8'h06;
        13'hAFB: rddata <= 8'h06;
        13'hAFC: rddata <= 8'h00;
        13'hAFD: rddata <= 8'h02;
        13'hAFE: rddata <= 8'h02;
        13'hAFF: rddata <= 8'h02;
        13'hB00: rddata <= 8'h00;
        13'hB01: rddata <= 8'h00;
        13'hB02: rddata <= 8'h00;
        13'hB03: rddata <= 8'h00;
        13'hB04: rddata <= 8'h00;
        13'hB05: rddata <= 8'h3C;
        13'hB06: rddata <= 8'h3C;
        13'hB07: rddata <= 8'h3C;
        13'hB08: rddata <= 8'h00;
        13'hB09: rddata <= 8'h0C;
        13'hB0A: rddata <= 8'h0C;
        13'hB0B: rddata <= 8'h0C;
        13'hB0C: rddata <= 8'h00;
        13'hB0D: rddata <= 8'h0C;
        13'hB0E: rddata <= 8'h0C;
        13'hB0F: rddata <= 8'h0C;
        13'hB10: rddata <= 8'h00;
        13'hB11: rddata <= 8'h0C;
        13'hB12: rddata <= 8'h0C;
        13'hB13: rddata <= 8'h0C;
        13'hB14: rddata <= 8'h00;
        13'hB15: rddata <= 8'h0C;
        13'hB16: rddata <= 8'h0C;
        13'hB17: rddata <= 8'h0C;
        13'hB18: rddata <= 8'h00;
        13'hB19: rddata <= 8'h0C;
        13'hB1A: rddata <= 8'h0C;
        13'hB1B: rddata <= 8'h0C;
        13'hB1C: rddata <= 8'h00;
        13'hB1D: rddata <= 8'h3C;
        13'hB1E: rddata <= 8'h3C;
        13'hB1F: rddata <= 8'h3C;
        13'hB20: rddata <= 8'h00;
        13'hB21: rddata <= 8'h00;
        13'hB22: rddata <= 8'h00;
        13'hB23: rddata <= 8'h00;
        13'hB24: rddata <= 8'h00;
        13'hB25: rddata <= 8'h18;
        13'hB26: rddata <= 8'h18;
        13'hB27: rddata <= 8'h18;
        13'hB28: rddata <= 8'h00;
        13'hB29: rddata <= 8'h3C;
        13'hB2A: rddata <= 8'h3C;
        13'hB2B: rddata <= 8'h3C;
        13'hB2C: rddata <= 8'h00;
        13'hB2D: rddata <= 8'h66;
        13'hB2E: rddata <= 8'h66;
        13'hB2F: rddata <= 8'h66;
        13'hB30: rddata <= 8'h00;
        13'hB31: rddata <= 8'h00;
        13'hB32: rddata <= 8'h00;
        13'hB33: rddata <= 8'h00;
        13'hB34: rddata <= 8'h00;
        13'hB35: rddata <= 8'h00;
        13'hB36: rddata <= 8'h00;
        13'hB37: rddata <= 8'h00;
        13'hB38: rddata <= 8'h00;
        13'hB39: rddata <= 8'h00;
        13'hB3A: rddata <= 8'h00;
        13'hB3B: rddata <= 8'h00;
        13'hB3C: rddata <= 8'h00;
        13'hB3D: rddata <= 8'h00;
        13'hB3E: rddata <= 8'h00;
        13'hB3F: rddata <= 8'h00;
        13'hB40: rddata <= 8'h00;
        13'hB41: rddata <= 8'h00;
        13'hB42: rddata <= 8'h00;
        13'hB43: rddata <= 8'h00;
        13'hB44: rddata <= 8'h00;
        13'hB45: rddata <= 8'h00;
        13'hB46: rddata <= 8'h00;
        13'hB47: rddata <= 8'h00;
        13'hB48: rddata <= 8'h00;
        13'hB49: rddata <= 8'h00;
        13'hB4A: rddata <= 8'h00;
        13'hB4B: rddata <= 8'h00;
        13'hB4C: rddata <= 8'h00;
        13'hB4D: rddata <= 8'h00;
        13'hB4E: rddata <= 8'h00;
        13'hB4F: rddata <= 8'h00;
        13'hB50: rddata <= 8'h00;
        13'hB51: rddata <= 8'h00;
        13'hB52: rddata <= 8'h00;
        13'hB53: rddata <= 8'h00;
        13'hB54: rddata <= 8'h00;
        13'hB55: rddata <= 8'h00;
        13'hB56: rddata <= 8'h00;
        13'hB57: rddata <= 8'h00;
        13'hB58: rddata <= 8'h00;
        13'hB59: rddata <= 8'h00;
        13'hB5A: rddata <= 8'h00;
        13'hB5B: rddata <= 8'h00;
        13'hB5C: rddata <= 8'h00;
        13'hB5D: rddata <= 8'h7E;
        13'hB5E: rddata <= 8'h7E;
        13'hB5F: rddata <= 8'h7E;
        13'hB60: rddata <= 8'h00;
        13'hB61: rddata <= 8'h00;
        13'hB62: rddata <= 8'h00;
        13'hB63: rddata <= 8'h00;
        13'hB64: rddata <= 8'h00;
        13'hB65: rddata <= 8'h18;
        13'hB66: rddata <= 8'h18;
        13'hB67: rddata <= 8'h18;
        13'hB68: rddata <= 8'h00;
        13'hB69: rddata <= 8'h18;
        13'hB6A: rddata <= 8'h18;
        13'hB6B: rddata <= 8'h18;
        13'hB6C: rddata <= 8'h00;
        13'hB6D: rddata <= 8'h0C;
        13'hB6E: rddata <= 8'h0C;
        13'hB6F: rddata <= 8'h0C;
        13'hB70: rddata <= 8'h00;
        13'hB71: rddata <= 8'h00;
        13'hB72: rddata <= 8'h00;
        13'hB73: rddata <= 8'h00;
        13'hB74: rddata <= 8'h00;
        13'hB75: rddata <= 8'h00;
        13'hB76: rddata <= 8'h00;
        13'hB77: rddata <= 8'h00;
        13'hB78: rddata <= 8'h00;
        13'hB79: rddata <= 8'h00;
        13'hB7A: rddata <= 8'h00;
        13'hB7B: rddata <= 8'h00;
        13'hB7C: rddata <= 8'h00;
        13'hB7D: rddata <= 8'h00;
        13'hB7E: rddata <= 8'h00;
        13'hB7F: rddata <= 8'h00;
        13'hB80: rddata <= 8'h00;
        13'hB81: rddata <= 8'h00;
        13'hB82: rddata <= 8'h00;
        13'hB83: rddata <= 8'h00;
        13'hB84: rddata <= 8'h00;
        13'hB85: rddata <= 8'h00;
        13'hB86: rddata <= 8'h00;
        13'hB87: rddata <= 8'h00;
        13'hB88: rddata <= 8'h00;
        13'hB89: rddata <= 8'h00;
        13'hB8A: rddata <= 8'h00;
        13'hB8B: rddata <= 8'h00;
        13'hB8C: rddata <= 8'h00;
        13'hB8D: rddata <= 8'h3C;
        13'hB8E: rddata <= 8'h3C;
        13'hB8F: rddata <= 8'h3C;
        13'hB90: rddata <= 8'h00;
        13'hB91: rddata <= 8'h06;
        13'hB92: rddata <= 8'h06;
        13'hB93: rddata <= 8'h06;
        13'hB94: rddata <= 8'h00;
        13'hB95: rddata <= 8'h3E;
        13'hB96: rddata <= 8'h3E;
        13'hB97: rddata <= 8'h3E;
        13'hB98: rddata <= 8'h00;
        13'hB99: rddata <= 8'h66;
        13'hB9A: rddata <= 8'h66;
        13'hB9B: rddata <= 8'h66;
        13'hB9C: rddata <= 8'h00;
        13'hB9D: rddata <= 8'h3E;
        13'hB9E: rddata <= 8'h3E;
        13'hB9F: rddata <= 8'h3E;
        13'hBA0: rddata <= 8'h00;
        13'hBA1: rddata <= 8'h00;
        13'hBA2: rddata <= 8'h00;
        13'hBA3: rddata <= 8'h00;
        13'hBA4: rddata <= 8'h00;
        13'hBA5: rddata <= 8'h60;
        13'hBA6: rddata <= 8'h60;
        13'hBA7: rddata <= 8'h60;
        13'hBA8: rddata <= 8'h00;
        13'hBA9: rddata <= 8'h60;
        13'hBAA: rddata <= 8'h60;
        13'hBAB: rddata <= 8'h60;
        13'hBAC: rddata <= 8'h00;
        13'hBAD: rddata <= 8'h7C;
        13'hBAE: rddata <= 8'h7C;
        13'hBAF: rddata <= 8'h7C;
        13'hBB0: rddata <= 8'h00;
        13'hBB1: rddata <= 8'h66;
        13'hBB2: rddata <= 8'h66;
        13'hBB3: rddata <= 8'h66;
        13'hBB4: rddata <= 8'h00;
        13'hBB5: rddata <= 8'h66;
        13'hBB6: rddata <= 8'h66;
        13'hBB7: rddata <= 8'h66;
        13'hBB8: rddata <= 8'h00;
        13'hBB9: rddata <= 8'h66;
        13'hBBA: rddata <= 8'h66;
        13'hBBB: rddata <= 8'h66;
        13'hBBC: rddata <= 8'h00;
        13'hBBD: rddata <= 8'h7C;
        13'hBBE: rddata <= 8'h7C;
        13'hBBF: rddata <= 8'h7C;
        13'hBC0: rddata <= 8'h00;
        13'hBC1: rddata <= 8'h00;
        13'hBC2: rddata <= 8'h00;
        13'hBC3: rddata <= 8'h00;
        13'hBC4: rddata <= 8'h00;
        13'hBC5: rddata <= 8'h00;
        13'hBC6: rddata <= 8'h00;
        13'hBC7: rddata <= 8'h00;
        13'hBC8: rddata <= 8'h00;
        13'hBC9: rddata <= 8'h00;
        13'hBCA: rddata <= 8'h00;
        13'hBCB: rddata <= 8'h00;
        13'hBCC: rddata <= 8'h00;
        13'hBCD: rddata <= 8'h3C;
        13'hBCE: rddata <= 8'h3C;
        13'hBCF: rddata <= 8'h3C;
        13'hBD0: rddata <= 8'h00;
        13'hBD1: rddata <= 8'h66;
        13'hBD2: rddata <= 8'h66;
        13'hBD3: rddata <= 8'h66;
        13'hBD4: rddata <= 8'h00;
        13'hBD5: rddata <= 8'h60;
        13'hBD6: rddata <= 8'h60;
        13'hBD7: rddata <= 8'h60;
        13'hBD8: rddata <= 8'h00;
        13'hBD9: rddata <= 8'h66;
        13'hBDA: rddata <= 8'h66;
        13'hBDB: rddata <= 8'h66;
        13'hBDC: rddata <= 8'h00;
        13'hBDD: rddata <= 8'h3C;
        13'hBDE: rddata <= 8'h3C;
        13'hBDF: rddata <= 8'h3C;
        13'hBE0: rddata <= 8'h00;
        13'hBE1: rddata <= 8'h00;
        13'hBE2: rddata <= 8'h00;
        13'hBE3: rddata <= 8'h00;
        13'hBE4: rddata <= 8'h00;
        13'hBE5: rddata <= 8'h06;
        13'hBE6: rddata <= 8'h06;
        13'hBE7: rddata <= 8'h06;
        13'hBE8: rddata <= 8'h00;
        13'hBE9: rddata <= 8'h06;
        13'hBEA: rddata <= 8'h06;
        13'hBEB: rddata <= 8'h06;
        13'hBEC: rddata <= 8'h00;
        13'hBED: rddata <= 8'h3E;
        13'hBEE: rddata <= 8'h3E;
        13'hBEF: rddata <= 8'h3E;
        13'hBF0: rddata <= 8'h00;
        13'hBF1: rddata <= 8'h66;
        13'hBF2: rddata <= 8'h66;
        13'hBF3: rddata <= 8'h66;
        13'hBF4: rddata <= 8'h00;
        13'hBF5: rddata <= 8'h66;
        13'hBF6: rddata <= 8'h66;
        13'hBF7: rddata <= 8'h66;
        13'hBF8: rddata <= 8'h00;
        13'hBF9: rddata <= 8'h66;
        13'hBFA: rddata <= 8'h66;
        13'hBFB: rddata <= 8'h66;
        13'hBFC: rddata <= 8'h00;
        13'hBFD: rddata <= 8'h3E;
        13'hBFE: rddata <= 8'h3E;
        13'hBFF: rddata <= 8'h3E;
        13'hC00: rddata <= 8'h00;
        13'hC01: rddata <= 8'h00;
        13'hC02: rddata <= 8'h00;
        13'hC03: rddata <= 8'h00;
        13'hC04: rddata <= 8'h00;
        13'hC05: rddata <= 8'h00;
        13'hC06: rddata <= 8'h00;
        13'hC07: rddata <= 8'h00;
        13'hC08: rddata <= 8'h00;
        13'hC09: rddata <= 8'h00;
        13'hC0A: rddata <= 8'h00;
        13'hC0B: rddata <= 8'h00;
        13'hC0C: rddata <= 8'h00;
        13'hC0D: rddata <= 8'h3C;
        13'hC0E: rddata <= 8'h3C;
        13'hC0F: rddata <= 8'h3C;
        13'hC10: rddata <= 8'h00;
        13'hC11: rddata <= 8'h66;
        13'hC12: rddata <= 8'h66;
        13'hC13: rddata <= 8'h66;
        13'hC14: rddata <= 8'h00;
        13'hC15: rddata <= 8'h7E;
        13'hC16: rddata <= 8'h7E;
        13'hC17: rddata <= 8'h7E;
        13'hC18: rddata <= 8'h00;
        13'hC19: rddata <= 8'h60;
        13'hC1A: rddata <= 8'h60;
        13'hC1B: rddata <= 8'h60;
        13'hC1C: rddata <= 8'h00;
        13'hC1D: rddata <= 8'h3C;
        13'hC1E: rddata <= 8'h3C;
        13'hC1F: rddata <= 8'h3C;
        13'hC20: rddata <= 8'h00;
        13'hC21: rddata <= 8'h00;
        13'hC22: rddata <= 8'h00;
        13'hC23: rddata <= 8'h00;
        13'hC24: rddata <= 8'h00;
        13'hC25: rddata <= 8'h3C;
        13'hC26: rddata <= 8'h3C;
        13'hC27: rddata <= 8'h3C;
        13'hC28: rddata <= 8'h00;
        13'hC29: rddata <= 8'h66;
        13'hC2A: rddata <= 8'h66;
        13'hC2B: rddata <= 8'h66;
        13'hC2C: rddata <= 8'h00;
        13'hC2D: rddata <= 8'h60;
        13'hC2E: rddata <= 8'h60;
        13'hC2F: rddata <= 8'h60;
        13'hC30: rddata <= 8'h00;
        13'hC31: rddata <= 8'hF8;
        13'hC32: rddata <= 8'hF8;
        13'hC33: rddata <= 8'hF8;
        13'hC34: rddata <= 8'h00;
        13'hC35: rddata <= 8'h60;
        13'hC36: rddata <= 8'h60;
        13'hC37: rddata <= 8'h60;
        13'hC38: rddata <= 8'h00;
        13'hC39: rddata <= 8'h60;
        13'hC3A: rddata <= 8'h60;
        13'hC3B: rddata <= 8'h60;
        13'hC3C: rddata <= 8'h00;
        13'hC3D: rddata <= 8'h60;
        13'hC3E: rddata <= 8'h60;
        13'hC3F: rddata <= 8'h60;
        13'hC40: rddata <= 8'h00;
        13'hC41: rddata <= 8'h00;
        13'hC42: rddata <= 8'h00;
        13'hC43: rddata <= 8'h00;
        13'hC44: rddata <= 8'h00;
        13'hC45: rddata <= 8'h00;
        13'hC46: rddata <= 8'h00;
        13'hC47: rddata <= 8'h00;
        13'hC48: rddata <= 8'h00;
        13'hC49: rddata <= 8'h00;
        13'hC4A: rddata <= 8'h00;
        13'hC4B: rddata <= 8'h00;
        13'hC4C: rddata <= 8'h00;
        13'hC4D: rddata <= 8'h3E;
        13'hC4E: rddata <= 8'h3E;
        13'hC4F: rddata <= 8'h3E;
        13'hC50: rddata <= 8'h00;
        13'hC51: rddata <= 8'h66;
        13'hC52: rddata <= 8'h66;
        13'hC53: rddata <= 8'h66;
        13'hC54: rddata <= 8'h00;
        13'hC55: rddata <= 8'h66;
        13'hC56: rddata <= 8'h66;
        13'hC57: rddata <= 8'h66;
        13'hC58: rddata <= 8'h00;
        13'hC59: rddata <= 8'h3E;
        13'hC5A: rddata <= 8'h3E;
        13'hC5B: rddata <= 8'h3E;
        13'hC5C: rddata <= 8'h00;
        13'hC5D: rddata <= 8'h06;
        13'hC5E: rddata <= 8'h06;
        13'hC5F: rddata <= 8'h06;
        13'hC60: rddata <= 8'h00;
        13'hC61: rddata <= 8'h3C;
        13'hC62: rddata <= 8'h3C;
        13'hC63: rddata <= 8'h3C;
        13'hC64: rddata <= 8'h00;
        13'hC65: rddata <= 8'h60;
        13'hC66: rddata <= 8'h60;
        13'hC67: rddata <= 8'h60;
        13'hC68: rddata <= 8'h00;
        13'hC69: rddata <= 8'h60;
        13'hC6A: rddata <= 8'h60;
        13'hC6B: rddata <= 8'h60;
        13'hC6C: rddata <= 8'h00;
        13'hC6D: rddata <= 8'h7C;
        13'hC6E: rddata <= 8'h7C;
        13'hC6F: rddata <= 8'h7C;
        13'hC70: rddata <= 8'h00;
        13'hC71: rddata <= 8'h66;
        13'hC72: rddata <= 8'h66;
        13'hC73: rddata <= 8'h66;
        13'hC74: rddata <= 8'h00;
        13'hC75: rddata <= 8'h66;
        13'hC76: rddata <= 8'h66;
        13'hC77: rddata <= 8'h66;
        13'hC78: rddata <= 8'h00;
        13'hC79: rddata <= 8'h66;
        13'hC7A: rddata <= 8'h66;
        13'hC7B: rddata <= 8'h66;
        13'hC7C: rddata <= 8'h00;
        13'hC7D: rddata <= 8'h66;
        13'hC7E: rddata <= 8'h66;
        13'hC7F: rddata <= 8'h66;
        13'hC80: rddata <= 8'h00;
        13'hC81: rddata <= 8'h00;
        13'hC82: rddata <= 8'h00;
        13'hC83: rddata <= 8'h00;
        13'hC84: rddata <= 8'h00;
        13'hC85: rddata <= 8'h18;
        13'hC86: rddata <= 8'h18;
        13'hC87: rddata <= 8'h18;
        13'hC88: rddata <= 8'h00;
        13'hC89: rddata <= 8'h00;
        13'hC8A: rddata <= 8'h00;
        13'hC8B: rddata <= 8'h00;
        13'hC8C: rddata <= 8'h00;
        13'hC8D: rddata <= 8'h18;
        13'hC8E: rddata <= 8'h18;
        13'hC8F: rddata <= 8'h18;
        13'hC90: rddata <= 8'h00;
        13'hC91: rddata <= 8'h18;
        13'hC92: rddata <= 8'h18;
        13'hC93: rddata <= 8'h18;
        13'hC94: rddata <= 8'h00;
        13'hC95: rddata <= 8'h18;
        13'hC96: rddata <= 8'h18;
        13'hC97: rddata <= 8'h18;
        13'hC98: rddata <= 8'h00;
        13'hC99: rddata <= 8'h18;
        13'hC9A: rddata <= 8'h18;
        13'hC9B: rddata <= 8'h18;
        13'hC9C: rddata <= 8'h00;
        13'hC9D: rddata <= 8'h0C;
        13'hC9E: rddata <= 8'h0C;
        13'hC9F: rddata <= 8'h0C;
        13'hCA0: rddata <= 8'h00;
        13'hCA1: rddata <= 8'h00;
        13'hCA2: rddata <= 8'h00;
        13'hCA3: rddata <= 8'h00;
        13'hCA4: rddata <= 8'h00;
        13'hCA5: rddata <= 8'h18;
        13'hCA6: rddata <= 8'h18;
        13'hCA7: rddata <= 8'h18;
        13'hCA8: rddata <= 8'h00;
        13'hCA9: rddata <= 8'h00;
        13'hCAA: rddata <= 8'h00;
        13'hCAB: rddata <= 8'h00;
        13'hCAC: rddata <= 8'h00;
        13'hCAD: rddata <= 8'h38;
        13'hCAE: rddata <= 8'h38;
        13'hCAF: rddata <= 8'h38;
        13'hCB0: rddata <= 8'h00;
        13'hCB1: rddata <= 8'h18;
        13'hCB2: rddata <= 8'h18;
        13'hCB3: rddata <= 8'h18;
        13'hCB4: rddata <= 8'h00;
        13'hCB5: rddata <= 8'h18;
        13'hCB6: rddata <= 8'h18;
        13'hCB7: rddata <= 8'h18;
        13'hCB8: rddata <= 8'h00;
        13'hCB9: rddata <= 8'h18;
        13'hCBA: rddata <= 8'h18;
        13'hCBB: rddata <= 8'h18;
        13'hCBC: rddata <= 8'h00;
        13'hCBD: rddata <= 8'h18;
        13'hCBE: rddata <= 8'h18;
        13'hCBF: rddata <= 8'h18;
        13'hCC0: rddata <= 8'h00;
        13'hCC1: rddata <= 8'h70;
        13'hCC2: rddata <= 8'h70;
        13'hCC3: rddata <= 8'h70;
        13'hCC4: rddata <= 8'h00;
        13'hCC5: rddata <= 8'h60;
        13'hCC6: rddata <= 8'h60;
        13'hCC7: rddata <= 8'h60;
        13'hCC8: rddata <= 8'h00;
        13'hCC9: rddata <= 8'h60;
        13'hCCA: rddata <= 8'h60;
        13'hCCB: rddata <= 8'h60;
        13'hCCC: rddata <= 8'h00;
        13'hCCD: rddata <= 8'h66;
        13'hCCE: rddata <= 8'h66;
        13'hCCF: rddata <= 8'h66;
        13'hCD0: rddata <= 8'h00;
        13'hCD1: rddata <= 8'h6C;
        13'hCD2: rddata <= 8'h6C;
        13'hCD3: rddata <= 8'h6C;
        13'hCD4: rddata <= 8'h00;
        13'hCD5: rddata <= 8'h78;
        13'hCD6: rddata <= 8'h78;
        13'hCD7: rddata <= 8'h78;
        13'hCD8: rddata <= 8'h00;
        13'hCD9: rddata <= 8'h6C;
        13'hCDA: rddata <= 8'h6C;
        13'hCDB: rddata <= 8'h6C;
        13'hCDC: rddata <= 8'h00;
        13'hCDD: rddata <= 8'h66;
        13'hCDE: rddata <= 8'h66;
        13'hCDF: rddata <= 8'h66;
        13'hCE0: rddata <= 8'h00;
        13'hCE1: rddata <= 8'h00;
        13'hCE2: rddata <= 8'h00;
        13'hCE3: rddata <= 8'h00;
        13'hCE4: rddata <= 8'h00;
        13'hCE5: rddata <= 8'h18;
        13'hCE6: rddata <= 8'h18;
        13'hCE7: rddata <= 8'h18;
        13'hCE8: rddata <= 8'h00;
        13'hCE9: rddata <= 8'h18;
        13'hCEA: rddata <= 8'h18;
        13'hCEB: rddata <= 8'h18;
        13'hCEC: rddata <= 8'h00;
        13'hCED: rddata <= 8'h18;
        13'hCEE: rddata <= 8'h18;
        13'hCEF: rddata <= 8'h18;
        13'hCF0: rddata <= 8'h00;
        13'hCF1: rddata <= 8'h18;
        13'hCF2: rddata <= 8'h18;
        13'hCF3: rddata <= 8'h18;
        13'hCF4: rddata <= 8'h00;
        13'hCF5: rddata <= 8'h18;
        13'hCF6: rddata <= 8'h18;
        13'hCF7: rddata <= 8'h18;
        13'hCF8: rddata <= 8'h00;
        13'hCF9: rddata <= 8'h18;
        13'hCFA: rddata <= 8'h18;
        13'hCFB: rddata <= 8'h18;
        13'hCFC: rddata <= 8'h00;
        13'hCFD: rddata <= 8'h0C;
        13'hCFE: rddata <= 8'h0C;
        13'hCFF: rddata <= 8'h0C;
        13'hD00: rddata <= 8'h00;
        13'hD01: rddata <= 8'h00;
        13'hD02: rddata <= 8'h00;
        13'hD03: rddata <= 8'h00;
        13'hD04: rddata <= 8'h00;
        13'hD05: rddata <= 8'h00;
        13'hD06: rddata <= 8'h00;
        13'hD07: rddata <= 8'h00;
        13'hD08: rddata <= 8'h00;
        13'hD09: rddata <= 8'h00;
        13'hD0A: rddata <= 8'h00;
        13'hD0B: rddata <= 8'h00;
        13'hD0C: rddata <= 8'h00;
        13'hD0D: rddata <= 8'hEC;
        13'hD0E: rddata <= 8'hEC;
        13'hD0F: rddata <= 8'hEC;
        13'hD10: rddata <= 8'h00;
        13'hD11: rddata <= 8'hFE;
        13'hD12: rddata <= 8'hFE;
        13'hD13: rddata <= 8'hFE;
        13'hD14: rddata <= 8'h00;
        13'hD15: rddata <= 8'hD6;
        13'hD16: rddata <= 8'hD6;
        13'hD17: rddata <= 8'hD6;
        13'hD18: rddata <= 8'h00;
        13'hD19: rddata <= 8'hD6;
        13'hD1A: rddata <= 8'hD6;
        13'hD1B: rddata <= 8'hD6;
        13'hD1C: rddata <= 8'h00;
        13'hD1D: rddata <= 8'hD6;
        13'hD1E: rddata <= 8'hD6;
        13'hD1F: rddata <= 8'hD6;
        13'hD20: rddata <= 8'h00;
        13'hD21: rddata <= 8'h00;
        13'hD22: rddata <= 8'h00;
        13'hD23: rddata <= 8'h00;
        13'hD24: rddata <= 8'h00;
        13'hD25: rddata <= 8'h00;
        13'hD26: rddata <= 8'h00;
        13'hD27: rddata <= 8'h00;
        13'hD28: rddata <= 8'h00;
        13'hD29: rddata <= 8'h00;
        13'hD2A: rddata <= 8'h00;
        13'hD2B: rddata <= 8'h00;
        13'hD2C: rddata <= 8'h00;
        13'hD2D: rddata <= 8'h7C;
        13'hD2E: rddata <= 8'h7C;
        13'hD2F: rddata <= 8'h7C;
        13'hD30: rddata <= 8'h00;
        13'hD31: rddata <= 8'h66;
        13'hD32: rddata <= 8'h66;
        13'hD33: rddata <= 8'h66;
        13'hD34: rddata <= 8'h00;
        13'hD35: rddata <= 8'h66;
        13'hD36: rddata <= 8'h66;
        13'hD37: rddata <= 8'h66;
        13'hD38: rddata <= 8'h00;
        13'hD39: rddata <= 8'h66;
        13'hD3A: rddata <= 8'h66;
        13'hD3B: rddata <= 8'h66;
        13'hD3C: rddata <= 8'h00;
        13'hD3D: rddata <= 8'h66;
        13'hD3E: rddata <= 8'h66;
        13'hD3F: rddata <= 8'h66;
        13'hD40: rddata <= 8'h00;
        13'hD41: rddata <= 8'h00;
        13'hD42: rddata <= 8'h00;
        13'hD43: rddata <= 8'h00;
        13'hD44: rddata <= 8'h00;
        13'hD45: rddata <= 8'h00;
        13'hD46: rddata <= 8'h00;
        13'hD47: rddata <= 8'h00;
        13'hD48: rddata <= 8'h00;
        13'hD49: rddata <= 8'h00;
        13'hD4A: rddata <= 8'h00;
        13'hD4B: rddata <= 8'h00;
        13'hD4C: rddata <= 8'h00;
        13'hD4D: rddata <= 8'h3C;
        13'hD4E: rddata <= 8'h3C;
        13'hD4F: rddata <= 8'h3C;
        13'hD50: rddata <= 8'h00;
        13'hD51: rddata <= 8'h66;
        13'hD52: rddata <= 8'h66;
        13'hD53: rddata <= 8'h66;
        13'hD54: rddata <= 8'h00;
        13'hD55: rddata <= 8'h66;
        13'hD56: rddata <= 8'h66;
        13'hD57: rddata <= 8'h66;
        13'hD58: rddata <= 8'h00;
        13'hD59: rddata <= 8'h66;
        13'hD5A: rddata <= 8'h66;
        13'hD5B: rddata <= 8'h66;
        13'hD5C: rddata <= 8'h00;
        13'hD5D: rddata <= 8'h3C;
        13'hD5E: rddata <= 8'h3C;
        13'hD5F: rddata <= 8'h3C;
        13'hD60: rddata <= 8'h00;
        13'hD61: rddata <= 8'h00;
        13'hD62: rddata <= 8'h00;
        13'hD63: rddata <= 8'h00;
        13'hD64: rddata <= 8'h00;
        13'hD65: rddata <= 8'h00;
        13'hD66: rddata <= 8'h00;
        13'hD67: rddata <= 8'h00;
        13'hD68: rddata <= 8'h00;
        13'hD69: rddata <= 8'h00;
        13'hD6A: rddata <= 8'h00;
        13'hD6B: rddata <= 8'h00;
        13'hD6C: rddata <= 8'h00;
        13'hD6D: rddata <= 8'h7C;
        13'hD6E: rddata <= 8'h7C;
        13'hD6F: rddata <= 8'h7C;
        13'hD70: rddata <= 8'h00;
        13'hD71: rddata <= 8'h66;
        13'hD72: rddata <= 8'h66;
        13'hD73: rddata <= 8'h66;
        13'hD74: rddata <= 8'h00;
        13'hD75: rddata <= 8'h66;
        13'hD76: rddata <= 8'h66;
        13'hD77: rddata <= 8'h66;
        13'hD78: rddata <= 8'h00;
        13'hD79: rddata <= 8'h7C;
        13'hD7A: rddata <= 8'h7C;
        13'hD7B: rddata <= 8'h7C;
        13'hD7C: rddata <= 8'h00;
        13'hD7D: rddata <= 8'h60;
        13'hD7E: rddata <= 8'h60;
        13'hD7F: rddata <= 8'h60;
        13'hD80: rddata <= 8'h00;
        13'hD81: rddata <= 8'h60;
        13'hD82: rddata <= 8'h60;
        13'hD83: rddata <= 8'h60;
        13'hD84: rddata <= 8'h00;
        13'hD85: rddata <= 8'h00;
        13'hD86: rddata <= 8'h00;
        13'hD87: rddata <= 8'h00;
        13'hD88: rddata <= 8'h00;
        13'hD89: rddata <= 8'h00;
        13'hD8A: rddata <= 8'h00;
        13'hD8B: rddata <= 8'h00;
        13'hD8C: rddata <= 8'h00;
        13'hD8D: rddata <= 8'h3E;
        13'hD8E: rddata <= 8'h3E;
        13'hD8F: rddata <= 8'h3E;
        13'hD90: rddata <= 8'h00;
        13'hD91: rddata <= 8'h66;
        13'hD92: rddata <= 8'h66;
        13'hD93: rddata <= 8'h66;
        13'hD94: rddata <= 8'h00;
        13'hD95: rddata <= 8'h66;
        13'hD96: rddata <= 8'h66;
        13'hD97: rddata <= 8'h66;
        13'hD98: rddata <= 8'h00;
        13'hD99: rddata <= 8'h3E;
        13'hD9A: rddata <= 8'h3E;
        13'hD9B: rddata <= 8'h3E;
        13'hD9C: rddata <= 8'h00;
        13'hD9D: rddata <= 8'h06;
        13'hD9E: rddata <= 8'h06;
        13'hD9F: rddata <= 8'h06;
        13'hDA0: rddata <= 8'h00;
        13'hDA1: rddata <= 8'h06;
        13'hDA2: rddata <= 8'h06;
        13'hDA3: rddata <= 8'h06;
        13'hDA4: rddata <= 8'h00;
        13'hDA5: rddata <= 8'h00;
        13'hDA6: rddata <= 8'h00;
        13'hDA7: rddata <= 8'h00;
        13'hDA8: rddata <= 8'h00;
        13'hDA9: rddata <= 8'h00;
        13'hDAA: rddata <= 8'h00;
        13'hDAB: rddata <= 8'h00;
        13'hDAC: rddata <= 8'h00;
        13'hDAD: rddata <= 8'h7C;
        13'hDAE: rddata <= 8'h7C;
        13'hDAF: rddata <= 8'h7C;
        13'hDB0: rddata <= 8'h00;
        13'hDB1: rddata <= 8'h66;
        13'hDB2: rddata <= 8'h66;
        13'hDB3: rddata <= 8'h66;
        13'hDB4: rddata <= 8'h00;
        13'hDB5: rddata <= 8'h60;
        13'hDB6: rddata <= 8'h60;
        13'hDB7: rddata <= 8'h60;
        13'hDB8: rddata <= 8'h00;
        13'hDB9: rddata <= 8'h60;
        13'hDBA: rddata <= 8'h60;
        13'hDBB: rddata <= 8'h60;
        13'hDBC: rddata <= 8'h00;
        13'hDBD: rddata <= 8'h60;
        13'hDBE: rddata <= 8'h60;
        13'hDBF: rddata <= 8'h60;
        13'hDC0: rddata <= 8'h00;
        13'hDC1: rddata <= 8'h00;
        13'hDC2: rddata <= 8'h00;
        13'hDC3: rddata <= 8'h00;
        13'hDC4: rddata <= 8'h00;
        13'hDC5: rddata <= 8'h00;
        13'hDC6: rddata <= 8'h00;
        13'hDC7: rddata <= 8'h00;
        13'hDC8: rddata <= 8'h00;
        13'hDC9: rddata <= 8'h00;
        13'hDCA: rddata <= 8'h00;
        13'hDCB: rddata <= 8'h00;
        13'hDCC: rddata <= 8'h00;
        13'hDCD: rddata <= 8'h3C;
        13'hDCE: rddata <= 8'h3C;
        13'hDCF: rddata <= 8'h3C;
        13'hDD0: rddata <= 8'h00;
        13'hDD1: rddata <= 8'h60;
        13'hDD2: rddata <= 8'h60;
        13'hDD3: rddata <= 8'h60;
        13'hDD4: rddata <= 8'h00;
        13'hDD5: rddata <= 8'h3C;
        13'hDD6: rddata <= 8'h3C;
        13'hDD7: rddata <= 8'h3C;
        13'hDD8: rddata <= 8'h00;
        13'hDD9: rddata <= 8'h06;
        13'hDDA: rddata <= 8'h06;
        13'hDDB: rddata <= 8'h06;
        13'hDDC: rddata <= 8'h00;
        13'hDDD: rddata <= 8'h3C;
        13'hDDE: rddata <= 8'h3C;
        13'hDDF: rddata <= 8'h3C;
        13'hDE0: rddata <= 8'h00;
        13'hDE1: rddata <= 8'h00;
        13'hDE2: rddata <= 8'h00;
        13'hDE3: rddata <= 8'h00;
        13'hDE4: rddata <= 8'h00;
        13'hDE5: rddata <= 8'h30;
        13'hDE6: rddata <= 8'h30;
        13'hDE7: rddata <= 8'h30;
        13'hDE8: rddata <= 8'h00;
        13'hDE9: rddata <= 8'h30;
        13'hDEA: rddata <= 8'h30;
        13'hDEB: rddata <= 8'h30;
        13'hDEC: rddata <= 8'h00;
        13'hDED: rddata <= 8'h7C;
        13'hDEE: rddata <= 8'h7C;
        13'hDEF: rddata <= 8'h7C;
        13'hDF0: rddata <= 8'h00;
        13'hDF1: rddata <= 8'h30;
        13'hDF2: rddata <= 8'h30;
        13'hDF3: rddata <= 8'h30;
        13'hDF4: rddata <= 8'h00;
        13'hDF5: rddata <= 8'h30;
        13'hDF6: rddata <= 8'h30;
        13'hDF7: rddata <= 8'h30;
        13'hDF8: rddata <= 8'h00;
        13'hDF9: rddata <= 8'h30;
        13'hDFA: rddata <= 8'h30;
        13'hDFB: rddata <= 8'h30;
        13'hDFC: rddata <= 8'h00;
        13'hDFD: rddata <= 8'h1C;
        13'hDFE: rddata <= 8'h1C;
        13'hDFF: rddata <= 8'h1C;
        13'hE00: rddata <= 8'h00;
        13'hE01: rddata <= 8'h00;
        13'hE02: rddata <= 8'h00;
        13'hE03: rddata <= 8'h00;
        13'hE04: rddata <= 8'h00;
        13'hE05: rddata <= 8'h00;
        13'hE06: rddata <= 8'h00;
        13'hE07: rddata <= 8'h00;
        13'hE08: rddata <= 8'h00;
        13'hE09: rddata <= 8'h00;
        13'hE0A: rddata <= 8'h00;
        13'hE0B: rddata <= 8'h00;
        13'hE0C: rddata <= 8'h00;
        13'hE0D: rddata <= 8'h66;
        13'hE0E: rddata <= 8'h66;
        13'hE0F: rddata <= 8'h66;
        13'hE10: rddata <= 8'h00;
        13'hE11: rddata <= 8'h66;
        13'hE12: rddata <= 8'h66;
        13'hE13: rddata <= 8'h66;
        13'hE14: rddata <= 8'h00;
        13'hE15: rddata <= 8'h66;
        13'hE16: rddata <= 8'h66;
        13'hE17: rddata <= 8'h66;
        13'hE18: rddata <= 8'h00;
        13'hE19: rddata <= 8'h66;
        13'hE1A: rddata <= 8'h66;
        13'hE1B: rddata <= 8'h66;
        13'hE1C: rddata <= 8'h00;
        13'hE1D: rddata <= 8'h3E;
        13'hE1E: rddata <= 8'h3E;
        13'hE1F: rddata <= 8'h3E;
        13'hE20: rddata <= 8'h00;
        13'hE21: rddata <= 8'h00;
        13'hE22: rddata <= 8'h00;
        13'hE23: rddata <= 8'h00;
        13'hE24: rddata <= 8'h00;
        13'hE25: rddata <= 8'h00;
        13'hE26: rddata <= 8'h00;
        13'hE27: rddata <= 8'h00;
        13'hE28: rddata <= 8'h00;
        13'hE29: rddata <= 8'h00;
        13'hE2A: rddata <= 8'h00;
        13'hE2B: rddata <= 8'h00;
        13'hE2C: rddata <= 8'h00;
        13'hE2D: rddata <= 8'h66;
        13'hE2E: rddata <= 8'h66;
        13'hE2F: rddata <= 8'h66;
        13'hE30: rddata <= 8'h00;
        13'hE31: rddata <= 8'h66;
        13'hE32: rddata <= 8'h66;
        13'hE33: rddata <= 8'h66;
        13'hE34: rddata <= 8'h00;
        13'hE35: rddata <= 8'h66;
        13'hE36: rddata <= 8'h66;
        13'hE37: rddata <= 8'h66;
        13'hE38: rddata <= 8'h00;
        13'hE39: rddata <= 8'h3C;
        13'hE3A: rddata <= 8'h3C;
        13'hE3B: rddata <= 8'h3C;
        13'hE3C: rddata <= 8'h00;
        13'hE3D: rddata <= 8'h18;
        13'hE3E: rddata <= 8'h18;
        13'hE3F: rddata <= 8'h18;
        13'hE40: rddata <= 8'h00;
        13'hE41: rddata <= 8'h00;
        13'hE42: rddata <= 8'h00;
        13'hE43: rddata <= 8'h00;
        13'hE44: rddata <= 8'h00;
        13'hE45: rddata <= 8'h00;
        13'hE46: rddata <= 8'h00;
        13'hE47: rddata <= 8'h00;
        13'hE48: rddata <= 8'h00;
        13'hE49: rddata <= 8'h00;
        13'hE4A: rddata <= 8'h00;
        13'hE4B: rddata <= 8'h00;
        13'hE4C: rddata <= 8'h00;
        13'hE4D: rddata <= 8'hC6;
        13'hE4E: rddata <= 8'hC6;
        13'hE4F: rddata <= 8'hC6;
        13'hE50: rddata <= 8'h00;
        13'hE51: rddata <= 8'hC6;
        13'hE52: rddata <= 8'hC6;
        13'hE53: rddata <= 8'hC6;
        13'hE54: rddata <= 8'h00;
        13'hE55: rddata <= 8'hD6;
        13'hE56: rddata <= 8'hD6;
        13'hE57: rddata <= 8'hD6;
        13'hE58: rddata <= 8'h00;
        13'hE59: rddata <= 8'hD6;
        13'hE5A: rddata <= 8'hD6;
        13'hE5B: rddata <= 8'hD6;
        13'hE5C: rddata <= 8'h00;
        13'hE5D: rddata <= 8'h6C;
        13'hE5E: rddata <= 8'h6C;
        13'hE5F: rddata <= 8'h6C;
        13'hE60: rddata <= 8'h00;
        13'hE61: rddata <= 8'h00;
        13'hE62: rddata <= 8'h00;
        13'hE63: rddata <= 8'h00;
        13'hE64: rddata <= 8'h00;
        13'hE65: rddata <= 8'h00;
        13'hE66: rddata <= 8'h00;
        13'hE67: rddata <= 8'h00;
        13'hE68: rddata <= 8'h00;
        13'hE69: rddata <= 8'h00;
        13'hE6A: rddata <= 8'h00;
        13'hE6B: rddata <= 8'h00;
        13'hE6C: rddata <= 8'h00;
        13'hE6D: rddata <= 8'h66;
        13'hE6E: rddata <= 8'h66;
        13'hE6F: rddata <= 8'h66;
        13'hE70: rddata <= 8'h00;
        13'hE71: rddata <= 8'h3C;
        13'hE72: rddata <= 8'h3C;
        13'hE73: rddata <= 8'h3C;
        13'hE74: rddata <= 8'h00;
        13'hE75: rddata <= 8'h18;
        13'hE76: rddata <= 8'h18;
        13'hE77: rddata <= 8'h18;
        13'hE78: rddata <= 8'h00;
        13'hE79: rddata <= 8'h3C;
        13'hE7A: rddata <= 8'h3C;
        13'hE7B: rddata <= 8'h3C;
        13'hE7C: rddata <= 8'h00;
        13'hE7D: rddata <= 8'h66;
        13'hE7E: rddata <= 8'h66;
        13'hE7F: rddata <= 8'h66;
        13'hE80: rddata <= 8'h00;
        13'hE81: rddata <= 8'h00;
        13'hE82: rddata <= 8'h00;
        13'hE83: rddata <= 8'h00;
        13'hE84: rddata <= 8'h00;
        13'hE85: rddata <= 8'h00;
        13'hE86: rddata <= 8'h00;
        13'hE87: rddata <= 8'h00;
        13'hE88: rddata <= 8'h00;
        13'hE89: rddata <= 8'h00;
        13'hE8A: rddata <= 8'h00;
        13'hE8B: rddata <= 8'h00;
        13'hE8C: rddata <= 8'h00;
        13'hE8D: rddata <= 8'h66;
        13'hE8E: rddata <= 8'h66;
        13'hE8F: rddata <= 8'h66;
        13'hE90: rddata <= 8'h00;
        13'hE91: rddata <= 8'h66;
        13'hE92: rddata <= 8'h66;
        13'hE93: rddata <= 8'h66;
        13'hE94: rddata <= 8'h00;
        13'hE95: rddata <= 8'h66;
        13'hE96: rddata <= 8'h66;
        13'hE97: rddata <= 8'h66;
        13'hE98: rddata <= 8'h00;
        13'hE99: rddata <= 8'h3E;
        13'hE9A: rddata <= 8'h3E;
        13'hE9B: rddata <= 8'h3E;
        13'hE9C: rddata <= 8'h00;
        13'hE9D: rddata <= 8'h06;
        13'hE9E: rddata <= 8'h06;
        13'hE9F: rddata <= 8'h06;
        13'hEA0: rddata <= 8'h00;
        13'hEA1: rddata <= 8'h3C;
        13'hEA2: rddata <= 8'h3C;
        13'hEA3: rddata <= 8'h3C;
        13'hEA4: rddata <= 8'h00;
        13'hEA5: rddata <= 8'h00;
        13'hEA6: rddata <= 8'h00;
        13'hEA7: rddata <= 8'h00;
        13'hEA8: rddata <= 8'h00;
        13'hEA9: rddata <= 8'h00;
        13'hEAA: rddata <= 8'h00;
        13'hEAB: rddata <= 8'h00;
        13'hEAC: rddata <= 8'h00;
        13'hEAD: rddata <= 8'h7E;
        13'hEAE: rddata <= 8'h7E;
        13'hEAF: rddata <= 8'h7E;
        13'hEB0: rddata <= 8'h00;
        13'hEB1: rddata <= 8'h0C;
        13'hEB2: rddata <= 8'h0C;
        13'hEB3: rddata <= 8'h0C;
        13'hEB4: rddata <= 8'h00;
        13'hEB5: rddata <= 8'h18;
        13'hEB6: rddata <= 8'h18;
        13'hEB7: rddata <= 8'h18;
        13'hEB8: rddata <= 8'h00;
        13'hEB9: rddata <= 8'h30;
        13'hEBA: rddata <= 8'h30;
        13'hEBB: rddata <= 8'h30;
        13'hEBC: rddata <= 8'h00;
        13'hEBD: rddata <= 8'h7E;
        13'hEBE: rddata <= 8'h7E;
        13'hEBF: rddata <= 8'h7E;
        13'hEC0: rddata <= 8'h00;
        13'hEC1: rddata <= 8'h00;
        13'hEC2: rddata <= 8'h00;
        13'hEC3: rddata <= 8'h00;
        13'hEC4: rddata <= 8'h00;
        13'hEC5: rddata <= 8'h0C;
        13'hEC6: rddata <= 8'h0C;
        13'hEC7: rddata <= 8'h0C;
        13'hEC8: rddata <= 8'h00;
        13'hEC9: rddata <= 8'h18;
        13'hECA: rddata <= 8'h18;
        13'hECB: rddata <= 8'h18;
        13'hECC: rddata <= 8'h00;
        13'hECD: rddata <= 8'h18;
        13'hECE: rddata <= 8'h18;
        13'hECF: rddata <= 8'h18;
        13'hED0: rddata <= 8'h00;
        13'hED1: rddata <= 8'h30;
        13'hED2: rddata <= 8'h30;
        13'hED3: rddata <= 8'h30;
        13'hED4: rddata <= 8'h00;
        13'hED5: rddata <= 8'h18;
        13'hED6: rddata <= 8'h18;
        13'hED7: rddata <= 8'h18;
        13'hED8: rddata <= 8'h00;
        13'hED9: rddata <= 8'h18;
        13'hEDA: rddata <= 8'h18;
        13'hEDB: rddata <= 8'h18;
        13'hEDC: rddata <= 8'h00;
        13'hEDD: rddata <= 8'h0C;
        13'hEDE: rddata <= 8'h0C;
        13'hEDF: rddata <= 8'h0C;
        13'hEE0: rddata <= 8'h00;
        13'hEE1: rddata <= 8'h00;
        13'hEE2: rddata <= 8'h00;
        13'hEE3: rddata <= 8'h00;
        13'hEE4: rddata <= 8'h00;
        13'hEE5: rddata <= 8'h18;
        13'hEE6: rddata <= 8'h18;
        13'hEE7: rddata <= 8'h18;
        13'hEE8: rddata <= 8'h00;
        13'hEE9: rddata <= 8'h18;
        13'hEEA: rddata <= 8'h18;
        13'hEEB: rddata <= 8'h18;
        13'hEEC: rddata <= 8'h00;
        13'hEED: rddata <= 8'h18;
        13'hEEE: rddata <= 8'h18;
        13'hEEF: rddata <= 8'h18;
        13'hEF0: rddata <= 8'h00;
        13'hEF1: rddata <= 8'h18;
        13'hEF2: rddata <= 8'h18;
        13'hEF3: rddata <= 8'h18;
        13'hEF4: rddata <= 8'h00;
        13'hEF5: rddata <= 8'h18;
        13'hEF6: rddata <= 8'h18;
        13'hEF7: rddata <= 8'h18;
        13'hEF8: rddata <= 8'h00;
        13'hEF9: rddata <= 8'h18;
        13'hEFA: rddata <= 8'h18;
        13'hEFB: rddata <= 8'h18;
        13'hEFC: rddata <= 8'h00;
        13'hEFD: rddata <= 8'h18;
        13'hEFE: rddata <= 8'h18;
        13'hEFF: rddata <= 8'h18;
        13'hF00: rddata <= 8'h00;
        13'hF01: rddata <= 8'h00;
        13'hF02: rddata <= 8'h00;
        13'hF03: rddata <= 8'h00;
        13'hF04: rddata <= 8'h00;
        13'hF05: rddata <= 8'h30;
        13'hF06: rddata <= 8'h30;
        13'hF07: rddata <= 8'h30;
        13'hF08: rddata <= 8'h00;
        13'hF09: rddata <= 8'h18;
        13'hF0A: rddata <= 8'h18;
        13'hF0B: rddata <= 8'h18;
        13'hF0C: rddata <= 8'h00;
        13'hF0D: rddata <= 8'h18;
        13'hF0E: rddata <= 8'h18;
        13'hF0F: rddata <= 8'h18;
        13'hF10: rddata <= 8'h00;
        13'hF11: rddata <= 8'h0C;
        13'hF12: rddata <= 8'h0C;
        13'hF13: rddata <= 8'h0C;
        13'hF14: rddata <= 8'h00;
        13'hF15: rddata <= 8'h18;
        13'hF16: rddata <= 8'h18;
        13'hF17: rddata <= 8'h18;
        13'hF18: rddata <= 8'h00;
        13'hF19: rddata <= 8'h18;
        13'hF1A: rddata <= 8'h18;
        13'hF1B: rddata <= 8'h18;
        13'hF1C: rddata <= 8'h00;
        13'hF1D: rddata <= 8'h30;
        13'hF1E: rddata <= 8'h30;
        13'hF1F: rddata <= 8'h30;
        13'hF20: rddata <= 8'h00;
        13'hF21: rddata <= 8'h00;
        13'hF22: rddata <= 8'h00;
        13'hF23: rddata <= 8'h00;
        13'hF24: rddata <= 8'h00;
        13'hF25: rddata <= 8'h00;
        13'hF26: rddata <= 8'h00;
        13'hF27: rddata <= 8'h00;
        13'hF28: rddata <= 8'h00;
        13'hF29: rddata <= 8'h00;
        13'hF2A: rddata <= 8'h00;
        13'hF2B: rddata <= 8'h00;
        13'hF2C: rddata <= 8'h00;
        13'hF2D: rddata <= 8'h00;
        13'hF2E: rddata <= 8'h00;
        13'hF2F: rddata <= 8'h00;
        13'hF30: rddata <= 8'h00;
        13'hF31: rddata <= 8'h3A;
        13'hF32: rddata <= 8'h3A;
        13'hF33: rddata <= 8'h3A;
        13'hF34: rddata <= 8'h00;
        13'hF35: rddata <= 8'h6E;
        13'hF36: rddata <= 8'h6E;
        13'hF37: rddata <= 8'h6E;
        13'hF38: rddata <= 8'h00;
        13'hF39: rddata <= 8'h00;
        13'hF3A: rddata <= 8'h00;
        13'hF3B: rddata <= 8'h00;
        13'hF3C: rddata <= 8'h00;
        13'hF3D: rddata <= 8'h00;
        13'hF3E: rddata <= 8'h00;
        13'hF3F: rddata <= 8'h00;
        13'hF40: rddata <= 8'h00;
        13'hF41: rddata <= 8'h00;
        13'hF42: rddata <= 8'h00;
        13'hF43: rddata <= 8'h00;
        13'hF44: rddata <= 8'h00;
        13'hF45: rddata <= 8'h3A;
        13'hF46: rddata <= 8'h07;
        13'hF47: rddata <= 8'hC0;
        13'hF48: rddata <= 8'h47;
        13'hF49: rddata <= 8'h3A;
        13'hF4A: rddata <= 8'h03;
        13'hF4B: rddata <= 8'hC0;
        13'hF4C: rddata <= 8'hB8;
        13'hF4D: rddata <= 8'h38;
        13'hF4E: rddata <= 8'h06;
        13'hF4F: rddata <= 8'h78;
        13'hF50: rddata <= 8'hD6;
        13'hF51: rddata <= 8'h01;
        13'hF52: rddata <= 8'h32;
        13'hF53: rddata <= 8'h03;
        13'hF54: rddata <= 8'hC0;
        13'hF55: rddata <= 8'hAF;
        13'hF56: rddata <= 8'hD3;
        13'hF57: rddata <= 8'hBF;
        13'hF58: rddata <= 8'h3E;
        13'hF59: rddata <= 8'h7F;
        13'hF5A: rddata <= 8'hD3;
        13'hF5B: rddata <= 8'hBF;
        13'hF5C: rddata <= 8'h3A;
        13'hF5D: rddata <= 8'h03;
        13'hF5E: rddata <= 8'hC0;
        13'hF5F: rddata <= 8'h87;
        13'hF60: rddata <= 8'h87;
        13'hF61: rddata <= 8'h87;
        13'hF62: rddata <= 8'hC6;
        13'hF63: rddata <= 8'h0E;
        13'hF64: rddata <= 8'hD3;
        13'hF65: rddata <= 8'hBE;
        13'hF66: rddata <= 8'h3E;
        13'hF67: rddata <= 8'hD0;
        13'hF68: rddata <= 8'hD3;
        13'hF69: rddata <= 8'hBE;
        13'hF6A: rddata <= 8'h3E;
        13'hF6B: rddata <= 8'h80;
        13'hF6C: rddata <= 8'hD3;
        13'hF6D: rddata <= 8'hBF;
        13'hF6E: rddata <= 8'h3E;
        13'hF6F: rddata <= 8'h7F;
        13'hF70: rddata <= 8'hD3;
        13'hF71: rddata <= 8'hBF;
        13'hF72: rddata <= 8'hAF;
        13'hF73: rddata <= 8'hD3;
        13'hF74: rddata <= 8'hBE;
        13'hF75: rddata <= 8'h3E;
        13'hF76: rddata <= 8'h1E;
        13'hF77: rddata <= 8'hD3;
        13'hF78: rddata <= 8'hBE;
        13'hF79: rddata <= 8'hC9;
        13'hF7A: rddata <= 8'hAF;
        13'hF7B: rddata <= 8'hD3;
        13'hF7C: rddata <= 8'hBF;
        13'hF7D: rddata <= 8'h3E;
        13'hF7E: rddata <= 8'h7F;
        13'hF7F: rddata <= 8'hD3;
        13'hF80: rddata <= 8'hBF;
        13'hF81: rddata <= 8'h3E;
        13'hF82: rddata <= 8'hD0;
        13'hF83: rddata <= 8'hD3;
        13'hF84: rddata <= 8'hBE;
        13'hF85: rddata <= 8'hC9;
        13'hF86: rddata <= 8'hAF;
        13'hF87: rddata <= 8'hD3;
        13'hF88: rddata <= 8'hBF;
        13'hF89: rddata <= 8'h3E;
        13'hF8A: rddata <= 8'h78;
        13'hF8B: rddata <= 8'hD3;
        13'hF8C: rddata <= 8'hBF;
        13'hF8D: rddata <= 8'hAF;
        13'hF8E: rddata <= 8'h0E;
        13'hF8F: rddata <= 8'h1C;
        13'hF90: rddata <= 8'h06;
        13'hF91: rddata <= 8'h20;
        13'hF92: rddata <= 8'hD3;
        13'hF93: rddata <= 8'hBE;
        13'hF94: rddata <= 8'hD3;
        13'hF95: rddata <= 8'hBE;
        13'hF96: rddata <= 8'h05;
        13'hF97: rddata <= 8'h20;
        13'hF98: rddata <= 8'hF9;
        13'hF99: rddata <= 8'h0D;
        13'hF9A: rddata <= 8'h20;
        13'hF9B: rddata <= 8'hF4;
        13'hF9C: rddata <= 8'hC9;
        13'hF9D: rddata <= 8'h26;
        13'hF9E: rddata <= 8'h00;
        13'hF9F: rddata <= 8'h3A;
        13'hFA0: rddata <= 8'h01;
        13'hFA1: rddata <= 8'hC0;
        13'hFA2: rddata <= 8'h6F;
        13'hFA3: rddata <= 8'h29;
        13'hFA4: rddata <= 8'h29;
        13'hFA5: rddata <= 8'h29;
        13'hFA6: rddata <= 8'h29;
        13'hFA7: rddata <= 8'h29;
        13'hFA8: rddata <= 8'h29;
        13'hFA9: rddata <= 8'h3A;
        13'hFAA: rddata <= 8'h00;
        13'hFAB: rddata <= 8'hC0;
        13'hFAC: rddata <= 8'h87;
        13'hFAD: rddata <= 8'h85;
        13'hFAE: rddata <= 8'hD3;
        13'hFAF: rddata <= 8'hBF;
        13'hFB0: rddata <= 8'h7C;
        13'hFB1: rddata <= 8'hC6;
        13'hFB2: rddata <= 8'h78;
        13'hFB3: rddata <= 8'hD3;
        13'hFB4: rddata <= 8'hBF;
        13'hFB5: rddata <= 8'hC9;
        13'hFB6: rddata <= 8'hFE;
        13'hFB7: rddata <= 8'h0A;
        13'hFB8: rddata <= 8'hCA;
        13'hFB9: rddata <= 8'hDD;
        13'hFBA: rddata <= 8'h0F;
        13'hFBB: rddata <= 8'hD6;
        13'hFBC: rddata <= 8'h20;
        13'hFBD: rddata <= 8'hFE;
        13'hFBE: rddata <= 8'h5F;
        13'hFBF: rddata <= 8'h38;
        13'hFC0: rddata <= 8'h01;
        13'hFC1: rddata <= 8'hAF;
        13'hFC2: rddata <= 8'hD3;
        13'hFC3: rddata <= 8'hBE;
        13'hFC4: rddata <= 8'hAF;
        13'hFC5: rddata <= 8'hD3;
        13'hFC6: rddata <= 8'hBE;
        13'hFC7: rddata <= 8'h3A;
        13'hFC8: rddata <= 8'h00;
        13'hFC9: rddata <= 8'hC0;
        13'hFCA: rddata <= 8'h3C;
        13'hFCB: rddata <= 8'h32;
        13'hFCC: rddata <= 8'h00;
        13'hFCD: rddata <= 8'hC0;
        13'hFCE: rddata <= 8'hFE;
        13'hFCF: rddata <= 8'h20;
        13'hFD0: rddata <= 8'hD8;
        13'hFD1: rddata <= 8'hAF;
        13'hFD2: rddata <= 8'h32;
        13'hFD3: rddata <= 8'h00;
        13'hFD4: rddata <= 8'hC0;
        13'hFD5: rddata <= 8'h3A;
        13'hFD6: rddata <= 8'h01;
        13'hFD7: rddata <= 8'hC0;
        13'hFD8: rddata <= 8'h3C;
        13'hFD9: rddata <= 8'h32;
        13'hFDA: rddata <= 8'h01;
        13'hFDB: rddata <= 8'hC0;
        13'hFDC: rddata <= 8'hC9;
        13'hFDD: rddata <= 8'hE5;
        13'hFDE: rddata <= 8'hAF;
        13'hFDF: rddata <= 8'h32;
        13'hFE0: rddata <= 8'h00;
        13'hFE1: rddata <= 8'hC0;
        13'hFE2: rddata <= 8'h3A;
        13'hFE3: rddata <= 8'h01;
        13'hFE4: rddata <= 8'hC0;
        13'hFE5: rddata <= 8'h3C;
        13'hFE6: rddata <= 8'h32;
        13'hFE7: rddata <= 8'h01;
        13'hFE8: rddata <= 8'hC0;
        13'hFE9: rddata <= 8'hCD;
        13'hFEA: rddata <= 8'h9D;
        13'hFEB: rddata <= 8'h0F;
        13'hFEC: rddata <= 8'hE1;
        13'hFED: rddata <= 8'hC9;
        13'hFEE: rddata <= 8'h7E;
        13'hFEF: rddata <= 8'hB7;
        13'hFF0: rddata <= 8'hC8;
        13'hFF1: rddata <= 8'hCD;
        13'hFF2: rddata <= 8'hB6;
        13'hFF3: rddata <= 8'h0F;
        13'hFF4: rddata <= 8'h23;
        13'hFF5: rddata <= 8'h18;
        13'hFF6: rddata <= 8'hF7;
        13'hFF7: rddata <= 8'hF5;
        13'hFF8: rddata <= 8'hDB;
        13'hFF9: rddata <= 8'h10;
        13'hFFA: rddata <= 8'hE6;
        13'hFFB: rddata <= 8'h01;
        13'hFFC: rddata <= 8'h28;
        13'hFFD: rddata <= 8'h04;
        13'hFFE: rddata <= 8'hDB;
        13'hFFF: rddata <= 8'h11;
        13'h1000: rddata <= 8'h18;
        13'h1001: rddata <= 8'hF6;
        13'h1002: rddata <= 8'h3E;
        13'h1003: rddata <= 8'h80;
        13'h1004: rddata <= 8'hD3;
        13'h1005: rddata <= 8'h10;
        13'h1006: rddata <= 8'hF1;
        13'h1007: rddata <= 8'hC3;
        13'h1008: rddata <= 8'h13;
        13'h1009: rddata <= 8'h10;
        13'h100A: rddata <= 8'hDB;
        13'h100B: rddata <= 8'h10;
        13'h100C: rddata <= 8'hE6;
        13'h100D: rddata <= 8'h01;
        13'h100E: rddata <= 8'h28;
        13'h100F: rddata <= 8'hFA;
        13'h1010: rddata <= 8'hDB;
        13'h1011: rddata <= 8'h11;
        13'h1012: rddata <= 8'hC9;
        13'h1013: rddata <= 8'hF5;
        13'h1014: rddata <= 8'hDB;
        13'h1015: rddata <= 8'h10;
        13'h1016: rddata <= 8'hE6;
        13'h1017: rddata <= 8'h02;
        13'h1018: rddata <= 8'h20;
        13'h1019: rddata <= 8'hFA;
        13'h101A: rddata <= 8'hF1;
        13'h101B: rddata <= 8'hD3;
        13'h101C: rddata <= 8'h11;
        13'h101D: rddata <= 8'hC9;
        13'h101E: rddata <= 8'h7E;
        13'h101F: rddata <= 8'hCD;
        13'h1020: rddata <= 8'h13;
        13'h1021: rddata <= 8'h10;
        13'h1022: rddata <= 8'hB7;
        13'h1023: rddata <= 8'hC8;
        13'h1024: rddata <= 8'h23;
        13'h1025: rddata <= 8'h18;
        13'h1026: rddata <= 8'hF7;
        13'h1027: rddata <= 8'h7A;
        13'h1028: rddata <= 8'hB3;
        13'h1029: rddata <= 8'hC8;
        13'h102A: rddata <= 8'hCD;
        13'h102B: rddata <= 8'h0A;
        13'h102C: rddata <= 8'h10;
        13'h102D: rddata <= 8'h77;
        13'h102E: rddata <= 8'h23;
        13'h102F: rddata <= 8'h1B;
        13'h1030: rddata <= 8'h18;
        13'h1031: rddata <= 8'hF5;
        13'h1032: rddata <= 8'h3E;
        13'h1033: rddata <= 8'h1F;
        13'h1034: rddata <= 8'hCD;
        13'h1035: rddata <= 8'hF7;
        13'h1036: rddata <= 8'h0F;
        13'h1037: rddata <= 8'hC3;
        13'h1038: rddata <= 8'h0A;
        13'h1039: rddata <= 8'h10;
        13'h103A: rddata <= 8'h3E;
        13'h103B: rddata <= 8'h16;
        13'h103C: rddata <= 8'hCD;
        13'h103D: rddata <= 8'hF7;
        13'h103E: rddata <= 8'h0F;
        13'h103F: rddata <= 8'hAF;
        13'h1040: rddata <= 8'hCD;
        13'h1041: rddata <= 8'h13;
        13'h1042: rddata <= 8'h10;
        13'h1043: rddata <= 8'hC3;
        13'h1044: rddata <= 8'h0A;
        13'h1045: rddata <= 8'h10;
        13'h1046: rddata <= 8'h3E;
        13'h1047: rddata <= 8'h18;
        13'h1048: rddata <= 8'hCD;
        13'h1049: rddata <= 8'hF7;
        13'h104A: rddata <= 8'h0F;
        13'h104B: rddata <= 8'hAF;
        13'h104C: rddata <= 8'hCD;
        13'h104D: rddata <= 8'h13;
        13'h104E: rddata <= 8'h10;
        13'h104F: rddata <= 8'hCD;
        13'h1050: rddata <= 8'h0A;
        13'h1051: rddata <= 8'h10;
        13'h1052: rddata <= 8'hB7;
        13'h1053: rddata <= 8'hC0;
        13'h1054: rddata <= 8'h21;
        13'h1055: rddata <= 8'h09;
        13'h1056: rddata <= 8'hC0;
        13'h1057: rddata <= 8'h11;
        13'h1058: rddata <= 8'h09;
        13'h1059: rddata <= 8'h00;
        13'h105A: rddata <= 8'hCD;
        13'h105B: rddata <= 8'h27;
        13'h105C: rddata <= 8'h10;
        13'h105D: rddata <= 8'h0E;
        13'h105E: rddata <= 8'h00;
        13'h105F: rddata <= 8'hCD;
        13'h1060: rddata <= 8'h0A;
        13'h1061: rddata <= 8'h10;
        13'h1062: rddata <= 8'h77;
        13'h1063: rddata <= 8'h23;
        13'h1064: rddata <= 8'hB7;
        13'h1065: rddata <= 8'h28;
        13'h1066: rddata <= 8'h03;
        13'h1067: rddata <= 8'h0C;
        13'h1068: rddata <= 8'h18;
        13'h1069: rddata <= 8'hF5;
        13'h106A: rddata <= 8'h79;
        13'h106B: rddata <= 8'h32;
        13'h106C: rddata <= 8'h08;
        13'h106D: rddata <= 8'hC0;
        13'h106E: rddata <= 8'h3A;
        13'h106F: rddata <= 8'h0D;
        13'h1070: rddata <= 8'hC0;
        13'h1071: rddata <= 8'hCB;
        13'h1072: rddata <= 8'h47;
        13'h1073: rddata <= 8'h20;
        13'h1074: rddata <= 8'h23;
        13'h1075: rddata <= 8'h3A;
        13'h1076: rddata <= 8'h08;
        13'h1077: rddata <= 8'hC0;
        13'h1078: rddata <= 8'hFE;
        13'h1079: rddata <= 8'h05;
        13'h107A: rddata <= 8'h38;
        13'h107B: rddata <= 8'hCA;
        13'h107C: rddata <= 8'hD6;
        13'h107D: rddata <= 8'h04;
        13'h107E: rddata <= 8'h32;
        13'h107F: rddata <= 8'h08;
        13'h1080: rddata <= 8'hC0;
        13'h1081: rddata <= 8'h21;
        13'h1082: rddata <= 8'h12;
        13'h1083: rddata <= 8'hC0;
        13'h1084: rddata <= 8'h06;
        13'h1085: rddata <= 8'h00;
        13'h1086: rddata <= 8'h4F;
        13'h1087: rddata <= 8'h09;
        13'h1088: rddata <= 8'hEB;
        13'h1089: rddata <= 8'h21;
        13'h108A: rddata <= 8'h9A;
        13'h108B: rddata <= 8'h10;
        13'h108C: rddata <= 8'h1A;
        13'h108D: rddata <= 8'hCD;
        13'h108E: rddata <= 8'h9F;
        13'h108F: rddata <= 8'h10;
        13'h1090: rddata <= 8'h13;
        13'h1091: rddata <= 8'hBE;
        13'h1092: rddata <= 8'h23;
        13'h1093: rddata <= 8'h20;
        13'h1094: rddata <= 8'hB1;
        13'h1095: rddata <= 8'hB7;
        13'h1096: rddata <= 8'h20;
        13'h1097: rddata <= 8'hF4;
        13'h1098: rddata <= 8'hAF;
        13'h1099: rddata <= 8'hC9;
        13'h109A: rddata <= 8'h2E;
        13'h109B: rddata <= 8'h53;
        13'h109C: rddata <= 8'h4D;
        13'h109D: rddata <= 8'h53;
        13'h109E: rddata <= 8'h00;
        13'h109F: rddata <= 8'hFE;
        13'h10A0: rddata <= 8'h61;
        13'h10A1: rddata <= 8'hD8;
        13'h10A2: rddata <= 8'hFE;
        13'h10A3: rddata <= 8'h7B;
        13'h10A4: rddata <= 8'hD0;
        13'h10A5: rddata <= 8'hD6;
        13'h10A6: rddata <= 8'h20;
        13'h10A7: rddata <= 8'hC9;
        13'h10A8: rddata <= 8'h3E;
        13'h10A9: rddata <= 8'h12;
        13'h10AA: rddata <= 8'hCD;
        13'h10AB: rddata <= 8'hF7;
        13'h10AC: rddata <= 8'h0F;
        13'h10AD: rddata <= 8'hAF;
        13'h10AE: rddata <= 8'hCD;
        13'h10AF: rddata <= 8'h13;
        13'h10B0: rddata <= 8'h10;
        13'h10B1: rddata <= 8'h7B;
        13'h10B2: rddata <= 8'hCD;
        13'h10B3: rddata <= 8'h13;
        13'h10B4: rddata <= 8'h10;
        13'h10B5: rddata <= 8'h7A;
        13'h10B6: rddata <= 8'hCD;
        13'h10B7: rddata <= 8'h13;
        13'h10B8: rddata <= 8'h10;
        13'h10B9: rddata <= 8'hCD;
        13'h10BA: rddata <= 8'h0A;
        13'h10BB: rddata <= 8'h10;
        13'h10BC: rddata <= 8'hCD;
        13'h10BD: rddata <= 8'h0A;
        13'h10BE: rddata <= 8'h10;
        13'h10BF: rddata <= 8'h5F;
        13'h10C0: rddata <= 8'hCD;
        13'h10C1: rddata <= 8'h0A;
        13'h10C2: rddata <= 8'h10;
        13'h10C3: rddata <= 8'h57;
        13'h10C4: rddata <= 8'hD5;
        13'h10C5: rddata <= 8'h7A;
        13'h10C6: rddata <= 8'hB3;
        13'h10C7: rddata <= 8'h28;
        13'h10C8: rddata <= 8'h08;
        13'h10C9: rddata <= 8'hCD;
        13'h10CA: rddata <= 8'h0A;
        13'h10CB: rddata <= 8'h10;
        13'h10CC: rddata <= 8'h77;
        13'h10CD: rddata <= 8'h23;
        13'h10CE: rddata <= 8'h1B;
        13'h10CF: rddata <= 8'h18;
        13'h10D0: rddata <= 8'hF4;
        13'h10D1: rddata <= 8'hD1;
        13'h10D2: rddata <= 8'hC9;
        13'h10D3: rddata <= 8'hAF;
        13'h10D4: rddata <= 8'h32;
        13'h10D5: rddata <= 8'hFD;
        13'h10D6: rddata <= 8'hFF;
        13'h10D7: rddata <= 8'h3C;
        13'h10D8: rddata <= 8'h32;
        13'h10D9: rddata <= 8'hFE;
        13'h10DA: rddata <= 8'hFF;
        13'h10DB: rddata <= 8'h3C;
        13'h10DC: rddata <= 8'h32;
        13'h10DD: rddata <= 8'hFF;
        13'h10DE: rddata <= 8'hFF;
        13'h10DF: rddata <= 8'hAF;
        13'h10E0: rddata <= 8'h32;
        13'h10E1: rddata <= 8'hFC;
        13'h10E2: rddata <= 8'hFF;
        13'h10E3: rddata <= 8'hC3;
        13'h10E4: rddata <= 8'h00;
        13'h10E5: rddata <= 8'h00;
        default:  rddata <= 8'h00;
    endcase

endmodule
