module rom(
    input  wire        clk,
    input  wire [13:0] addr,
    output reg   [7:0] rddata);

    always @(posedge clk)
        case (addr)
            14'h0000: rddata <= 8'hC3; 14'h0001: rddata <= 8'h00; 14'h0002: rddata <= 8'h20; 14'h0003: rddata <= 8'h82;
            14'h0004: rddata <= 8'h06; 14'h0005: rddata <= 8'h22; 14'h0006: rddata <= 8'h0B; 14'h0007: rddata <= 8'h00;
            14'h0008: rddata <= 8'h7E; 14'h0009: rddata <= 8'hE3; 14'h000A: rddata <= 8'hBE; 14'h000B: rddata <= 8'h23;
            14'h000C: rddata <= 8'hE3; 14'h000D: rddata <= 8'hC2; 14'h000E: rddata <= 8'hC4; 14'h000F: rddata <= 8'h03;
            14'h0010: rddata <= 8'h23; 14'h0011: rddata <= 8'h7E; 14'h0012: rddata <= 8'hFE; 14'h0013: rddata <= 8'h3A;
            14'h0014: rddata <= 8'hD0; 14'h0015: rddata <= 8'hC3; 14'h0016: rddata <= 8'h70; 14'h0017: rddata <= 8'h06;
            14'h0018: rddata <= 8'hC3; 14'h0019: rddata <= 8'h8A; 14'h001A: rddata <= 8'h19; 14'h001B: rddata <= 8'h00;
            14'h001C: rddata <= 8'h00; 14'h001D: rddata <= 8'h00; 14'h001E: rddata <= 8'h00; 14'h001F: rddata <= 8'h00;
            14'h0020: rddata <= 8'h7C; 14'h0021: rddata <= 8'h92; 14'h0022: rddata <= 8'hC0; 14'h0023: rddata <= 8'h7D;
            14'h0024: rddata <= 8'h93; 14'h0025: rddata <= 8'hC9; 14'h0026: rddata <= 8'h00; 14'h0027: rddata <= 8'h00;
            14'h0028: rddata <= 8'h3A; 14'h0029: rddata <= 8'hE7; 14'h002A: rddata <= 8'h38; 14'h002B: rddata <= 8'hB7;
            14'h002C: rddata <= 8'hC2; 14'h002D: rddata <= 8'hEB; 14'h002E: rddata <= 8'h14; 14'h002F: rddata <= 8'hC9;
            14'h0030: rddata <= 8'hDD; 14'h0031: rddata <= 8'h2A; 14'h0032: rddata <= 8'h06; 14'h0033: rddata <= 8'h38;
            14'h0034: rddata <= 8'hDD; 14'h0035: rddata <= 8'hE9; 14'h0036: rddata <= 8'h00; 14'h0037: rddata <= 8'h00;
            14'h0038: rddata <= 8'hC3; 14'h0039: rddata <= 8'h03; 14'h003A: rddata <= 8'h38; 14'h003B: rddata <= 8'hD9;
            14'h003C: rddata <= 8'hE1; 14'h003D: rddata <= 8'h23; 14'h003E: rddata <= 8'hE5; 14'h003F: rddata <= 8'hD9;
            14'h0040: rddata <= 8'hC9; 14'h0041: rddata <= 8'h31; 14'h0042: rddata <= 8'hA0; 14'h0043: rddata <= 8'h38;
            14'h0044: rddata <= 8'h3E; 14'h0045: rddata <= 8'h0B; 14'h0046: rddata <= 8'hCD; 14'h0047: rddata <= 8'h94;
            14'h0048: rddata <= 8'h1D; 14'h0049: rddata <= 8'h2A; 14'h004A: rddata <= 8'h01; 14'h004B: rddata <= 8'h38;
            14'h004C: rddata <= 8'h36; 14'h004D: rddata <= 8'h20; 14'h004E: rddata <= 8'h3E; 14'h004F: rddata <= 8'h07;
            14'h0050: rddata <= 8'hCD; 14'h0051: rddata <= 8'h94; 14'h0052: rddata <= 8'h1D; 14'h0053: rddata <= 8'hAF;
            14'h0054: rddata <= 8'hD3; 14'h0055: rddata <= 8'hFF; 14'h0056: rddata <= 8'h21; 14'h0057: rddata <= 8'hFF;
            14'h0058: rddata <= 8'h2F; 14'h0059: rddata <= 8'h22; 14'h005A: rddata <= 8'h5D; 14'h005B: rddata <= 8'h38;
            14'h005C: rddata <= 8'h11; 14'h005D: rddata <= 8'h11; 14'h005E: rddata <= 8'hE0; 14'h005F: rddata <= 8'h21;
            14'h0060: rddata <= 8'h81; 14'h0061: rddata <= 8'h00; 14'h0062: rddata <= 8'h1B; 14'h0063: rddata <= 8'h1B;
            14'h0064: rddata <= 8'h23; 14'h0065: rddata <= 8'h1A; 14'h0066: rddata <= 8'h0F; 14'h0067: rddata <= 8'h0F;
            14'h0068: rddata <= 8'h83; 14'h0069: rddata <= 8'hBE; 14'h006A: rddata <= 8'h28; 14'h006B: rddata <= 8'hF6;
            14'h006C: rddata <= 8'h7E; 14'h006D: rddata <= 8'hB7; 14'h006E: rddata <= 8'h20; 14'h006F: rddata <= 8'h19;
            14'h0070: rddata <= 8'hEB; 14'h0071: rddata <= 8'h06; 14'h0072: rddata <= 8'h0C; 14'h0073: rddata <= 8'h86;
            14'h0074: rddata <= 8'h23; 14'h0075: rddata <= 8'h80; 14'h0076: rddata <= 8'h05; 14'h0077: rddata <= 8'h20;
            14'h0078: rddata <= 8'hFA; 14'h0079: rddata <= 8'hAE; 14'h007A: rddata <= 8'hD3; 14'h007B: rddata <= 8'hFF;
            14'h007C: rddata <= 8'h32; 14'h007D: rddata <= 8'h09; 14'h007E: rddata <= 8'h38; 14'h007F: rddata <= 8'hC3;
            14'h0080: rddata <= 8'h06; 14'h0081: rddata <= 8'h20; 14'h0082: rddata <= 8'h2B; 14'h0083: rddata <= 8'h37;
            14'h0084: rddata <= 8'h24; 14'h0085: rddata <= 8'h24; 14'h0086: rddata <= 8'h33; 14'h0087: rddata <= 8'h2C;
            14'h0088: rddata <= 8'h00; 14'h0089: rddata <= 8'h11; 14'h008A: rddata <= 8'hA1; 14'h008B: rddata <= 8'h31;
            14'h008C: rddata <= 8'h21; 14'h008D: rddata <= 8'hB0; 14'h008E: rddata <= 8'h00; 14'h008F: rddata <= 8'h01;
            14'h0090: rddata <= 8'h05; 14'h0091: rddata <= 8'h00; 14'h0092: rddata <= 8'hED; 14'h0093: rddata <= 8'hB0;
            14'h0094: rddata <= 8'h11; 14'h0095: rddata <= 8'h10; 14'h0096: rddata <= 8'h32; 14'h0097: rddata <= 8'h21;
            14'h0098: rddata <= 8'hB5; 14'h0099: rddata <= 8'h00; 14'h009A: rddata <= 8'h01; 14'h009B: rddata <= 8'h19;
            14'h009C: rddata <= 8'h00; 14'h009D: rddata <= 8'hED; 14'h009E: rddata <= 8'hB0; 14'h009F: rddata <= 8'h06;
            14'h00A0: rddata <= 8'h03; 14'h00A1: rddata <= 8'hCD; 14'h00A2: rddata <= 8'hCF; 14'h00A3: rddata <= 8'h00;
            14'h00A4: rddata <= 8'h06; 14'h00A5: rddata <= 8'h02; 14'h00A6: rddata <= 8'hCD; 14'h00A7: rddata <= 8'hCF;
            14'h00A8: rddata <= 8'h00; 14'h00A9: rddata <= 8'h06; 14'h00AA: rddata <= 8'h06; 14'h00AB: rddata <= 8'hCD;
            14'h00AC: rddata <= 8'hCF; 14'h00AD: rddata <= 8'h00; 14'h00AE: rddata <= 8'h18; 14'h00AF: rddata <= 8'hEF;
            14'h00B0: rddata <= 8'h42; 14'h00B1: rddata <= 8'h41; 14'h00B2: rddata <= 8'h53; 14'h00B3: rddata <= 8'h49;
            14'h00B4: rddata <= 8'h43; 14'h00B5: rddata <= 8'h50; 14'h00B6: rddata <= 8'h72; 14'h00B7: rddata <= 8'h65;
            14'h00B8: rddata <= 8'h73; 14'h00B9: rddata <= 8'h73; 14'h00BA: rddata <= 8'h20; 14'h00BB: rddata <= 8'h52;
            14'h00BC: rddata <= 8'h45; 14'h00BD: rddata <= 8'h54; 14'h00BE: rddata <= 8'h55; 14'h00BF: rddata <= 8'h52;
            14'h00C0: rddata <= 8'h4E; 14'h00C1: rddata <= 8'h20; 14'h00C2: rddata <= 8'h6B; 14'h00C3: rddata <= 8'h65;
            14'h00C4: rddata <= 8'h79; 14'h00C5: rddata <= 8'h20; 14'h00C6: rddata <= 8'h74; 14'h00C7: rddata <= 8'h6F;
            14'h00C8: rddata <= 8'h20; 14'h00C9: rddata <= 8'h73; 14'h00CA: rddata <= 8'h74; 14'h00CB: rddata <= 8'h61;
            14'h00CC: rddata <= 8'h72; 14'h00CD: rddata <= 8'h74; 14'h00CE: rddata <= 8'h00; 14'h00CF: rddata <= 8'h21;
            14'h00D0: rddata <= 8'h00; 14'h00D1: rddata <= 8'h34; 14'h00D2: rddata <= 8'h70; 14'h00D3: rddata <= 8'h23;
            14'h00D4: rddata <= 8'h7C; 14'h00D5: rddata <= 8'hFE; 14'h00D6: rddata <= 8'h38; 14'h00D7: rddata <= 8'h20;
            14'h00D8: rddata <= 8'hF9; 14'h00D9: rddata <= 8'h21; 14'h00DA: rddata <= 8'h00; 14'h00DB: rddata <= 8'h40;
            14'h00DC: rddata <= 8'hCD; 14'h00DD: rddata <= 8'h80; 14'h00DE: rddata <= 8'h1E; 14'h00DF: rddata <= 8'hFE;
            14'h00E0: rddata <= 8'h0D; 14'h00E1: rddata <= 8'h28; 14'h00E2: rddata <= 8'h1A; 14'h00E3: rddata <= 8'hFE;
            14'h00E4: rddata <= 8'h03; 14'h00E5: rddata <= 8'h28; 14'h00E6: rddata <= 8'h06; 14'h00E7: rddata <= 8'h2B;
            14'h00E8: rddata <= 8'h7C; 14'h00E9: rddata <= 8'hB5; 14'h00EA: rddata <= 8'h20; 14'h00EB: rddata <= 8'hF0;
            14'h00EC: rddata <= 8'hC9; 14'h00ED: rddata <= 8'h3E; 14'h00EE: rddata <= 8'h0B; 14'h00EF: rddata <= 8'hCD;
            14'h00F0: rddata <= 8'h72; 14'h00F1: rddata <= 8'h1D; 14'h00F2: rddata <= 8'h3A; 14'h00F3: rddata <= 8'h09;
            14'h00F4: rddata <= 8'h38; 14'h00F5: rddata <= 8'hD3; 14'h00F6: rddata <= 8'hFF; 14'h00F7: rddata <= 8'hCD;
            14'h00F8: rddata <= 8'hE5; 14'h00F9: rddata <= 8'h0B; 14'h00FA: rddata <= 8'hCD; 14'h00FB: rddata <= 8'h40;
            14'h00FC: rddata <= 8'h1A; 14'h00FD: rddata <= 8'h21; 14'h00FE: rddata <= 8'h87; 14'h00FF: rddata <= 8'h01;
            14'h0100: rddata <= 8'h01; 14'h0101: rddata <= 8'h51; 14'h0102: rddata <= 8'h00; 14'h0103: rddata <= 8'h11;
            14'h0104: rddata <= 8'h03; 14'h0105: rddata <= 8'h38; 14'h0106: rddata <= 8'hED; 14'h0107: rddata <= 8'hB0;
            14'h0108: rddata <= 8'hAF; 14'h0109: rddata <= 8'h32; 14'h010A: rddata <= 8'hA9; 14'h010B: rddata <= 8'h38;
            14'h010C: rddata <= 8'h32; 14'h010D: rddata <= 8'h00; 14'h010E: rddata <= 8'h39; 14'h010F: rddata <= 8'hC3;
            14'h0110: rddata <= 8'h03; 14'h0111: rddata <= 8'h20; 14'h0112: rddata <= 8'h23; 14'h0113: rddata <= 8'h4E;
            14'h0114: rddata <= 8'h7C; 14'h0115: rddata <= 8'hB5; 14'h0116: rddata <= 8'h28; 14'h0117: rddata <= 8'h0B;
            14'h0118: rddata <= 8'hA9; 14'h0119: rddata <= 8'h77; 14'h011A: rddata <= 8'h46; 14'h011B: rddata <= 8'h2F;
            14'h011C: rddata <= 8'h77; 14'h011D: rddata <= 8'h7E; 14'h011E: rddata <= 8'h2F; 14'h011F: rddata <= 8'h71;
            14'h0120: rddata <= 8'hB8; 14'h0121: rddata <= 8'h28; 14'h0122: rddata <= 8'hEF; 14'h0123: rddata <= 8'h2B;
            14'h0124: rddata <= 8'h11; 14'h0125: rddata <= 8'h2C; 14'h0126: rddata <= 8'h3A; 14'h0127: rddata <= 8'hE7;
            14'h0128: rddata <= 8'hDA; 14'h0129: rddata <= 8'hB7; 14'h012A: rddata <= 8'h0B; 14'h012B: rddata <= 8'h11;
            14'h012C: rddata <= 8'hCE; 14'h012D: rddata <= 8'hFF; 14'h012E: rddata <= 8'h22; 14'h012F: rddata <= 8'hAD;
            14'h0130: rddata <= 8'h38; 14'h0131: rddata <= 8'h19; 14'h0132: rddata <= 8'h22; 14'h0133: rddata <= 8'h4B;
            14'h0134: rddata <= 8'h38; 14'h0135: rddata <= 8'hCD; 14'h0136: rddata <= 8'hBE; 14'h0137: rddata <= 8'h0B;
            14'h0138: rddata <= 8'hCD; 14'h0139: rddata <= 8'hF2; 14'h013A: rddata <= 8'h1F; 14'h013B: rddata <= 8'h31;
            14'h013C: rddata <= 8'h65; 14'h013D: rddata <= 8'h38; 14'h013E: rddata <= 8'hCD; 14'h013F: rddata <= 8'hE5;
            14'h0140: rddata <= 8'h0B; 14'h0141: rddata <= 8'h21; 14'h0142: rddata <= 8'h05; 14'h0143: rddata <= 8'h20;
            14'h0144: rddata <= 8'h11; 14'h0145: rddata <= 8'h82; 14'h0146: rddata <= 8'h00; 14'h0147: rddata <= 8'h1A;
            14'h0148: rddata <= 8'hB7; 14'h0149: rddata <= 8'hCA; 14'h014A: rddata <= 8'hE8; 14'h014B: rddata <= 8'h1F;
            14'h014C: rddata <= 8'hBE; 14'h014D: rddata <= 8'h20; 14'h014E: rddata <= 8'h04; 14'h014F: rddata <= 8'h2B;
            14'h0150: rddata <= 8'h13; 14'h0151: rddata <= 8'h18; 14'h0152: rddata <= 8'hF4; 14'h0153: rddata <= 8'hED;
            14'h0154: rddata <= 8'h5F; 14'h0155: rddata <= 8'h17; 14'h0156: rddata <= 8'hAF; 14'h0157: rddata <= 8'hD3;
            14'h0158: rddata <= 8'hFF; 14'h0159: rddata <= 8'h32; 14'h015A: rddata <= 8'h09; 14'h015B: rddata <= 8'h38;
            14'h015C: rddata <= 8'hC3; 14'h015D: rddata <= 8'h02; 14'h015E: rddata <= 8'h04; 14'h015F: rddata <= 8'h0B;
            14'h0160: rddata <= 8'h43; 14'h0161: rddata <= 8'h6F; 14'h0162: rddata <= 8'h70; 14'h0163: rddata <= 8'h79;
            14'h0164: rddata <= 8'h72; 14'h0165: rddata <= 8'h69; 14'h0166: rddata <= 8'h67; 14'h0167: rddata <= 8'h68;
            14'h0168: rddata <= 8'h74; 14'h0169: rddata <= 8'h20; 14'h016A: rddata <= 8'h05; 14'h016B: rddata <= 8'h20;
            14'h016C: rddata <= 8'h31; 14'h016D: rddata <= 8'h39; 14'h016E: rddata <= 8'h38; 14'h016F: rddata <= 8'h32;
            14'h0170: rddata <= 8'h20; 14'h0171: rddata <= 8'h62; 14'h0172: rddata <= 8'h79; 14'h0173: rddata <= 8'h20;
            14'h0174: rddata <= 8'h4D; 14'h0175: rddata <= 8'h69; 14'h0176: rddata <= 8'h63; 14'h0177: rddata <= 8'h72;
            14'h0178: rddata <= 8'h6F; 14'h0179: rddata <= 8'h73; 14'h017A: rddata <= 8'h6F; 14'h017B: rddata <= 8'h66;
            14'h017C: rddata <= 8'h74; 14'h017D: rddata <= 8'h20; 14'h017E: rddata <= 8'h49; 14'h017F: rddata <= 8'h6E;
            14'h0180: rddata <= 8'h63; 14'h0181: rddata <= 8'h2E; 14'h0182: rddata <= 8'h20; 14'h0183: rddata <= 8'h53;
            14'h0184: rddata <= 8'h32; 14'h0185: rddata <= 8'h0A; 14'h0186: rddata <= 8'h00; 14'h0187: rddata <= 8'hC3;
            14'h0188: rddata <= 8'h97; 14'h0189: rddata <= 8'h06; 14'h018A: rddata <= 8'h3B; 14'h018B: rddata <= 8'h00;
            14'h018C: rddata <= 8'h00; 14'h018D: rddata <= 8'hA3; 14'h018E: rddata <= 8'h00; 14'h018F: rddata <= 8'h00;
            14'h0190: rddata <= 8'h00; 14'h0191: rddata <= 8'h20; 14'h0192: rddata <= 8'h00; 14'h0193: rddata <= 8'h00;
            14'h0194: rddata <= 8'hD6; 14'h0195: rddata <= 8'h00; 14'h0196: rddata <= 8'h6F; 14'h0197: rddata <= 8'h7C;
            14'h0198: rddata <= 8'hDE; 14'h0199: rddata <= 8'h00; 14'h019A: rddata <= 8'h67; 14'h019B: rddata <= 8'h78;
            14'h019C: rddata <= 8'hDE; 14'h019D: rddata <= 8'h00; 14'h019E: rddata <= 8'h47; 14'h019F: rddata <= 8'h3E;
            14'h01A0: rddata <= 8'h00; 14'h01A1: rddata <= 8'hC9; 14'h01A2: rddata <= 8'h00; 14'h01A3: rddata <= 8'h00;
            14'h01A4: rddata <= 8'h00; 14'h01A5: rddata <= 8'h35; 14'h01A6: rddata <= 8'h4A; 14'h01A7: rddata <= 8'hCA;
            14'h01A8: rddata <= 8'h99; 14'h01A9: rddata <= 8'h39; 14'h01AA: rddata <= 8'h1C; 14'h01AB: rddata <= 8'h76;
            14'h01AC: rddata <= 8'h98; 14'h01AD: rddata <= 8'h22; 14'h01AE: rddata <= 8'h95; 14'h01AF: rddata <= 8'hB3;
            14'h01B0: rddata <= 8'h98; 14'h01B1: rddata <= 8'h0A; 14'h01B2: rddata <= 8'hDD; 14'h01B3: rddata <= 8'h47;
            14'h01B4: rddata <= 8'h98; 14'h01B5: rddata <= 8'h53; 14'h01B6: rddata <= 8'hD1; 14'h01B7: rddata <= 8'h99;
            14'h01B8: rddata <= 8'h99; 14'h01B9: rddata <= 8'h0A; 14'h01BA: rddata <= 8'h1A; 14'h01BB: rddata <= 8'h9F;
            14'h01BC: rddata <= 8'h98; 14'h01BD: rddata <= 8'h65; 14'h01BE: rddata <= 8'hBC; 14'h01BF: rddata <= 8'hCD;
            14'h01C0: rddata <= 8'h98; 14'h01C1: rddata <= 8'hD6; 14'h01C2: rddata <= 8'h77; 14'h01C3: rddata <= 8'h3E;
            14'h01C4: rddata <= 8'h98; 14'h01C5: rddata <= 8'h52; 14'h01C6: rddata <= 8'hC7; 14'h01C7: rddata <= 8'h4F;
            14'h01C8: rddata <= 8'h80; 14'h01C9: rddata <= 8'h00; 14'h01CA: rddata <= 8'h00; 14'h01CB: rddata <= 8'h00;
            14'h01CC: rddata <= 8'h28; 14'h01CD: rddata <= 8'h0E; 14'h01CE: rddata <= 8'h00; 14'h01CF: rddata <= 8'h64;
            14'h01D0: rddata <= 8'h39; 14'h01D1: rddata <= 8'hFE; 14'h01D2: rddata <= 8'hFF; 14'h01D3: rddata <= 8'h01;
            14'h01D4: rddata <= 8'h39; 14'h01D5: rddata <= 8'h21; 14'h01D6: rddata <= 8'h0C; 14'h01D7: rddata <= 8'hBC;
            14'h01D8: rddata <= 8'h05; 14'h01D9: rddata <= 8'h13; 14'h01DA: rddata <= 8'h0D; 14'h01DB: rddata <= 8'h1C;
            14'h01DC: rddata <= 8'h07; 14'h01DD: rddata <= 8'h93; 14'h01DE: rddata <= 8'h08; 14'h01DF: rddata <= 8'hCC;
            14'h01E0: rddata <= 8'h10; 14'h01E1: rddata <= 8'hBE; 14'h01E2: rddata <= 8'h08; 14'h01E3: rddata <= 8'h31;
            14'h01E4: rddata <= 8'h07; 14'h01E5: rddata <= 8'hDC; 14'h01E6: rddata <= 8'h06; 14'h01E7: rddata <= 8'hBE;
            14'h01E8: rddata <= 8'h06; 14'h01E9: rddata <= 8'h9C; 14'h01EA: rddata <= 8'h07; 14'h01EB: rddata <= 8'h05;
            14'h01EC: rddata <= 8'h0C; 14'h01ED: rddata <= 8'hCB; 14'h01EE: rddata <= 8'h06; 14'h01EF: rddata <= 8'hF8;
            14'h01F0: rddata <= 8'h06; 14'h01F1: rddata <= 8'h1E; 14'h01F2: rddata <= 8'h07; 14'h01F3: rddata <= 8'h1F;
            14'h01F4: rddata <= 8'h0C; 14'h01F5: rddata <= 8'h80; 14'h01F6: rddata <= 8'h07; 14'h01F7: rddata <= 8'hB5;
            14'h01F8: rddata <= 8'h07; 14'h01F9: rddata <= 8'h15; 14'h01FA: rddata <= 8'h1B; 14'h01FB: rddata <= 8'h3B;
            14'h01FC: rddata <= 8'h0B; 14'h01FD: rddata <= 8'h6D; 14'h01FE: rddata <= 8'h0B; 14'h01FF: rddata <= 8'hBC;
            14'h0200: rddata <= 8'h07; 14'h0201: rddata <= 8'h4B; 14'h0202: rddata <= 8'h0C; 14'h0203: rddata <= 8'h6C;
            14'h0204: rddata <= 8'h05; 14'h0205: rddata <= 8'h67; 14'h0206: rddata <= 8'h05; 14'h0207: rddata <= 8'hCD;
            14'h0208: rddata <= 8'h0C; 14'h0209: rddata <= 8'h2C; 14'h020A: rddata <= 8'h1C; 14'h020B: rddata <= 8'h08;
            14'h020C: rddata <= 8'h1C; 14'h020D: rddata <= 8'h4F; 14'h020E: rddata <= 8'h1A; 14'h020F: rddata <= 8'h4C;
            14'h0210: rddata <= 8'h1A; 14'h0211: rddata <= 8'hD6; 14'h0212: rddata <= 8'h1A; 14'h0213: rddata <= 8'hBD;
            14'h0214: rddata <= 8'h0B; 14'h0215: rddata <= 8'hF5; 14'h0216: rddata <= 8'h14; 14'h0217: rddata <= 8'hB1;
            14'h0218: rddata <= 8'h15; 14'h0219: rddata <= 8'h09; 14'h021A: rddata <= 8'h15; 14'h021B: rddata <= 8'h03;
            14'h021C: rddata <= 8'h38; 14'h021D: rddata <= 8'hA8; 14'h021E: rddata <= 8'h10; 14'h021F: rddata <= 8'h2E;
            14'h0220: rddata <= 8'h0B; 14'h0221: rddata <= 8'h33; 14'h0222: rddata <= 8'h0B; 14'h0223: rddata <= 8'h75;
            14'h0224: rddata <= 8'h17; 14'h0225: rddata <= 8'h66; 14'h0226: rddata <= 8'h18; 14'h0227: rddata <= 8'h85;
            14'h0228: rddata <= 8'h13; 14'h0229: rddata <= 8'hCD; 14'h022A: rddata <= 8'h17; 14'h022B: rddata <= 8'hD7;
            14'h022C: rddata <= 8'h18; 14'h022D: rddata <= 8'hDD; 14'h022E: rddata <= 8'h18; 14'h022F: rddata <= 8'h70;
            14'h0230: rddata <= 8'h19; 14'h0231: rddata <= 8'h85; 14'h0232: rddata <= 8'h19; 14'h0233: rddata <= 8'h63;
            14'h0234: rddata <= 8'h0B; 14'h0235: rddata <= 8'hF3; 14'h0236: rddata <= 8'h0F; 14'h0237: rddata <= 8'h29;
            14'h0238: rddata <= 8'h0E; 14'h0239: rddata <= 8'h84; 14'h023A: rddata <= 8'h10; 14'h023B: rddata <= 8'h02;
            14'h023C: rddata <= 8'h10; 14'h023D: rddata <= 8'h13; 14'h023E: rddata <= 8'h10; 14'h023F: rddata <= 8'h21;
            14'h0240: rddata <= 8'h10; 14'h0241: rddata <= 8'h50; 14'h0242: rddata <= 8'h10; 14'h0243: rddata <= 8'h59;
            14'h0244: rddata <= 8'h10; 14'h0245: rddata <= 8'hC5; 14'h0246: rddata <= 8'h4E; 14'h0247: rddata <= 8'h44;
            14'h0248: rddata <= 8'hC6; 14'h0249: rddata <= 8'h4F; 14'h024A: rddata <= 8'h52; 14'h024B: rddata <= 8'hCE;
            14'h024C: rddata <= 8'h45; 14'h024D: rddata <= 8'h58; 14'h024E: rddata <= 8'h54; 14'h024F: rddata <= 8'hC4;
            14'h0250: rddata <= 8'h41; 14'h0251: rddata <= 8'h54; 14'h0252: rddata <= 8'h41; 14'h0253: rddata <= 8'hC9;
            14'h0254: rddata <= 8'h4E; 14'h0255: rddata <= 8'h50; 14'h0256: rddata <= 8'h55; 14'h0257: rddata <= 8'h54;
            14'h0258: rddata <= 8'hC4; 14'h0259: rddata <= 8'h49; 14'h025A: rddata <= 8'h4D; 14'h025B: rddata <= 8'hD2;
            14'h025C: rddata <= 8'h45; 14'h025D: rddata <= 8'h41; 14'h025E: rddata <= 8'h44; 14'h025F: rddata <= 8'hCC;
            14'h0260: rddata <= 8'h45; 14'h0261: rddata <= 8'h54; 14'h0262: rddata <= 8'hC7; 14'h0263: rddata <= 8'h4F;
            14'h0264: rddata <= 8'h54; 14'h0265: rddata <= 8'h4F; 14'h0266: rddata <= 8'hD2; 14'h0267: rddata <= 8'h55;
            14'h0268: rddata <= 8'h4E; 14'h0269: rddata <= 8'hC9; 14'h026A: rddata <= 8'h46; 14'h026B: rddata <= 8'hD2;
            14'h026C: rddata <= 8'h45; 14'h026D: rddata <= 8'h53; 14'h026E: rddata <= 8'h54; 14'h026F: rddata <= 8'h4F;
            14'h0270: rddata <= 8'h52; 14'h0271: rddata <= 8'h45; 14'h0272: rddata <= 8'hC7; 14'h0273: rddata <= 8'h4F;
            14'h0274: rddata <= 8'h53; 14'h0275: rddata <= 8'h55; 14'h0276: rddata <= 8'h42; 14'h0277: rddata <= 8'hD2;
            14'h0278: rddata <= 8'h45; 14'h0279: rddata <= 8'h54; 14'h027A: rddata <= 8'h55; 14'h027B: rddata <= 8'h52;
            14'h027C: rddata <= 8'h4E; 14'h027D: rddata <= 8'hD2; 14'h027E: rddata <= 8'h45; 14'h027F: rddata <= 8'h4D;
            14'h0280: rddata <= 8'hD3; 14'h0281: rddata <= 8'h54; 14'h0282: rddata <= 8'h4F; 14'h0283: rddata <= 8'h50;
            14'h0284: rddata <= 8'hCF; 14'h0285: rddata <= 8'h4E; 14'h0286: rddata <= 8'hCC; 14'h0287: rddata <= 8'h50;
            14'h0288: rddata <= 8'h52; 14'h0289: rddata <= 8'h49; 14'h028A: rddata <= 8'h4E; 14'h028B: rddata <= 8'h54;
            14'h028C: rddata <= 8'hC3; 14'h028D: rddata <= 8'h4F; 14'h028E: rddata <= 8'h50; 14'h028F: rddata <= 8'h59;
            14'h0290: rddata <= 8'hC4; 14'h0291: rddata <= 8'h45; 14'h0292: rddata <= 8'h46; 14'h0293: rddata <= 8'hD0;
            14'h0294: rddata <= 8'h4F; 14'h0295: rddata <= 8'h4B; 14'h0296: rddata <= 8'h45; 14'h0297: rddata <= 8'hD0;
            14'h0298: rddata <= 8'h52; 14'h0299: rddata <= 8'h49; 14'h029A: rddata <= 8'h4E; 14'h029B: rddata <= 8'h54;
            14'h029C: rddata <= 8'hC3; 14'h029D: rddata <= 8'h4F; 14'h029E: rddata <= 8'h4E; 14'h029F: rddata <= 8'h54;
            14'h02A0: rddata <= 8'hCC; 14'h02A1: rddata <= 8'h49; 14'h02A2: rddata <= 8'h53; 14'h02A3: rddata <= 8'h54;
            14'h02A4: rddata <= 8'hCC; 14'h02A5: rddata <= 8'h4C; 14'h02A6: rddata <= 8'h49; 14'h02A7: rddata <= 8'h53;
            14'h02A8: rddata <= 8'h54; 14'h02A9: rddata <= 8'hC3; 14'h02AA: rddata <= 8'h4C; 14'h02AB: rddata <= 8'h45;
            14'h02AC: rddata <= 8'h41; 14'h02AD: rddata <= 8'h52; 14'h02AE: rddata <= 8'hC3; 14'h02AF: rddata <= 8'h4C;
            14'h02B0: rddata <= 8'h4F; 14'h02B1: rddata <= 8'h41; 14'h02B2: rddata <= 8'h44; 14'h02B3: rddata <= 8'hC3;
            14'h02B4: rddata <= 8'h53; 14'h02B5: rddata <= 8'h41; 14'h02B6: rddata <= 8'h56; 14'h02B7: rddata <= 8'h45;
            14'h02B8: rddata <= 8'hD0; 14'h02B9: rddata <= 8'h53; 14'h02BA: rddata <= 8'h45; 14'h02BB: rddata <= 8'h54;
            14'h02BC: rddata <= 8'hD0; 14'h02BD: rddata <= 8'h52; 14'h02BE: rddata <= 8'h45; 14'h02BF: rddata <= 8'h53;
            14'h02C0: rddata <= 8'h45; 14'h02C1: rddata <= 8'h54; 14'h02C2: rddata <= 8'hD3; 14'h02C3: rddata <= 8'h4F;
            14'h02C4: rddata <= 8'h55; 14'h02C5: rddata <= 8'h4E; 14'h02C6: rddata <= 8'h44; 14'h02C7: rddata <= 8'hCE;
            14'h02C8: rddata <= 8'h45; 14'h02C9: rddata <= 8'h57; 14'h02CA: rddata <= 8'hD4; 14'h02CB: rddata <= 8'h41;
            14'h02CC: rddata <= 8'h42; 14'h02CD: rddata <= 8'h28; 14'h02CE: rddata <= 8'hD4; 14'h02CF: rddata <= 8'h4F;
            14'h02D0: rddata <= 8'hC6; 14'h02D1: rddata <= 8'h4E; 14'h02D2: rddata <= 8'hD3; 14'h02D3: rddata <= 8'h50;
            14'h02D4: rddata <= 8'h43; 14'h02D5: rddata <= 8'h28; 14'h02D6: rddata <= 8'hC9; 14'h02D7: rddata <= 8'h4E;
            14'h02D8: rddata <= 8'h4B; 14'h02D9: rddata <= 8'h45; 14'h02DA: rddata <= 8'h59; 14'h02DB: rddata <= 8'h24;
            14'h02DC: rddata <= 8'hD4; 14'h02DD: rddata <= 8'h48; 14'h02DE: rddata <= 8'h45; 14'h02DF: rddata <= 8'h4E;
            14'h02E0: rddata <= 8'hCE; 14'h02E1: rddata <= 8'h4F; 14'h02E2: rddata <= 8'h54; 14'h02E3: rddata <= 8'hD3;
            14'h02E4: rddata <= 8'h54; 14'h02E5: rddata <= 8'h45; 14'h02E6: rddata <= 8'h50; 14'h02E7: rddata <= 8'hAB;
            14'h02E8: rddata <= 8'hAD; 14'h02E9: rddata <= 8'hAA; 14'h02EA: rddata <= 8'hAF; 14'h02EB: rddata <= 8'hDE;
            14'h02EC: rddata <= 8'hC1; 14'h02ED: rddata <= 8'h4E; 14'h02EE: rddata <= 8'h44; 14'h02EF: rddata <= 8'hCF;
            14'h02F0: rddata <= 8'h52; 14'h02F1: rddata <= 8'hBE; 14'h02F2: rddata <= 8'hBD; 14'h02F3: rddata <= 8'hBC;
            14'h02F4: rddata <= 8'hD3; 14'h02F5: rddata <= 8'h47; 14'h02F6: rddata <= 8'h4E; 14'h02F7: rddata <= 8'hC9;
            14'h02F8: rddata <= 8'h4E; 14'h02F9: rddata <= 8'h54; 14'h02FA: rddata <= 8'hC1; 14'h02FB: rddata <= 8'h42;
            14'h02FC: rddata <= 8'h53; 14'h02FD: rddata <= 8'hD5; 14'h02FE: rddata <= 8'h53; 14'h02FF: rddata <= 8'h52;
            14'h0300: rddata <= 8'hC6; 14'h0301: rddata <= 8'h52; 14'h0302: rddata <= 8'h45; 14'h0303: rddata <= 8'hCC;
            14'h0304: rddata <= 8'h50; 14'h0305: rddata <= 8'h4F; 14'h0306: rddata <= 8'h53; 14'h0307: rddata <= 8'hD0;
            14'h0308: rddata <= 8'h4F; 14'h0309: rddata <= 8'h53; 14'h030A: rddata <= 8'hD3; 14'h030B: rddata <= 8'h51;
            14'h030C: rddata <= 8'h52; 14'h030D: rddata <= 8'hD2; 14'h030E: rddata <= 8'h4E; 14'h030F: rddata <= 8'h44;
            14'h0310: rddata <= 8'hCC; 14'h0311: rddata <= 8'h4F; 14'h0312: rddata <= 8'h47; 14'h0313: rddata <= 8'hC5;
            14'h0314: rddata <= 8'h58; 14'h0315: rddata <= 8'h50; 14'h0316: rddata <= 8'hC3; 14'h0317: rddata <= 8'h4F;
            14'h0318: rddata <= 8'h53; 14'h0319: rddata <= 8'hD3; 14'h031A: rddata <= 8'h49; 14'h031B: rddata <= 8'h4E;
            14'h031C: rddata <= 8'hD4; 14'h031D: rddata <= 8'h41; 14'h031E: rddata <= 8'h4E; 14'h031F: rddata <= 8'hC1;
            14'h0320: rddata <= 8'h54; 14'h0321: rddata <= 8'h4E; 14'h0322: rddata <= 8'hD0; 14'h0323: rddata <= 8'h45;
            14'h0324: rddata <= 8'h45; 14'h0325: rddata <= 8'h4B; 14'h0326: rddata <= 8'hCC; 14'h0327: rddata <= 8'h45;
            14'h0328: rddata <= 8'h4E; 14'h0329: rddata <= 8'hD3; 14'h032A: rddata <= 8'h54; 14'h032B: rddata <= 8'h52;
            14'h032C: rddata <= 8'h24; 14'h032D: rddata <= 8'hD6; 14'h032E: rddata <= 8'h41; 14'h032F: rddata <= 8'h4C;
            14'h0330: rddata <= 8'hC1; 14'h0331: rddata <= 8'h53; 14'h0332: rddata <= 8'h43; 14'h0333: rddata <= 8'hC3;
            14'h0334: rddata <= 8'h48; 14'h0335: rddata <= 8'h52; 14'h0336: rddata <= 8'h24; 14'h0337: rddata <= 8'hCC;
            14'h0338: rddata <= 8'h45; 14'h0339: rddata <= 8'h46; 14'h033A: rddata <= 8'h54; 14'h033B: rddata <= 8'h24;
            14'h033C: rddata <= 8'hD2; 14'h033D: rddata <= 8'h49; 14'h033E: rddata <= 8'h47; 14'h033F: rddata <= 8'h48;
            14'h0340: rddata <= 8'h54; 14'h0341: rddata <= 8'h24; 14'h0342: rddata <= 8'hCD; 14'h0343: rddata <= 8'h49;
            14'h0344: rddata <= 8'h44; 14'h0345: rddata <= 8'h24; 14'h0346: rddata <= 8'hD0; 14'h0347: rddata <= 8'h4F;
            14'h0348: rddata <= 8'h49; 14'h0349: rddata <= 8'h4E; 14'h034A: rddata <= 8'h54; 14'h034B: rddata <= 8'h80;
            14'h034C: rddata <= 8'h79; 14'h034D: rddata <= 8'h5C; 14'h034E: rddata <= 8'h16; 14'h034F: rddata <= 8'h79;
            14'h0350: rddata <= 8'h5C; 14'h0351: rddata <= 8'h12; 14'h0352: rddata <= 8'h7C; 14'h0353: rddata <= 8'hC9;
            14'h0354: rddata <= 8'h13; 14'h0355: rddata <= 8'h7C; 14'h0356: rddata <= 8'h2D; 14'h0357: rddata <= 8'h14;
            14'h0358: rddata <= 8'h7F; 14'h0359: rddata <= 8'h7E; 14'h035A: rddata <= 8'h17; 14'h035B: rddata <= 8'h50;
            14'h035C: rddata <= 8'hA9; 14'h035D: rddata <= 8'h0A; 14'h035E: rddata <= 8'h46; 14'h035F: rddata <= 8'hA8;
            14'h0360: rddata <= 8'h0A; 14'h0361: rddata <= 8'h20; 14'h0362: rddata <= 8'h45; 14'h0363: rddata <= 8'h72;
            14'h0364: rddata <= 8'h72; 14'h0365: rddata <= 8'h6F; 14'h0366: rddata <= 8'h72; 14'h0367: rddata <= 8'h07;
            14'h0368: rddata <= 8'h00; 14'h0369: rddata <= 8'h20; 14'h036A: rddata <= 8'h69; 14'h036B: rddata <= 8'h6E;
            14'h036C: rddata <= 8'h20; 14'h036D: rddata <= 8'h00; 14'h036E: rddata <= 8'h4F; 14'h036F: rddata <= 8'h6B;
            14'h0370: rddata <= 8'h0D; 14'h0371: rddata <= 8'h0A; 14'h0372: rddata <= 8'h00; 14'h0373: rddata <= 8'h42;
            14'h0374: rddata <= 8'h72; 14'h0375: rddata <= 8'h65; 14'h0376: rddata <= 8'h61; 14'h0377: rddata <= 8'h6B;
            14'h0378: rddata <= 8'h00; 14'h0379: rddata <= 8'h4E; 14'h037A: rddata <= 8'h46; 14'h037B: rddata <= 8'h53;
            14'h037C: rddata <= 8'h4E; 14'h037D: rddata <= 8'h52; 14'h037E: rddata <= 8'h47; 14'h037F: rddata <= 8'h4F;
            14'h0380: rddata <= 8'h44; 14'h0381: rddata <= 8'h46; 14'h0382: rddata <= 8'h43; 14'h0383: rddata <= 8'h4F;
            14'h0384: rddata <= 8'h56; 14'h0385: rddata <= 8'h4F; 14'h0386: rddata <= 8'h4D; 14'h0387: rddata <= 8'h55;
            14'h0388: rddata <= 8'h4C; 14'h0389: rddata <= 8'h42; 14'h038A: rddata <= 8'h53; 14'h038B: rddata <= 8'h44;
            14'h038C: rddata <= 8'h44; 14'h038D: rddata <= 8'h2F; 14'h038E: rddata <= 8'h30; 14'h038F: rddata <= 8'h49;
            14'h0390: rddata <= 8'h44; 14'h0391: rddata <= 8'h54; 14'h0392: rddata <= 8'h4D; 14'h0393: rddata <= 8'h4F;
            14'h0394: rddata <= 8'h53; 14'h0395: rddata <= 8'h4C; 14'h0396: rddata <= 8'h53; 14'h0397: rddata <= 8'h53;
            14'h0398: rddata <= 8'h54; 14'h0399: rddata <= 8'h43; 14'h039A: rddata <= 8'h4E; 14'h039B: rddata <= 8'h55;
            14'h039C: rddata <= 8'h46; 14'h039D: rddata <= 8'h4D; 14'h039E: rddata <= 8'h4F; 14'h039F: rddata <= 8'h21;
            14'h03A0: rddata <= 8'h04; 14'h03A1: rddata <= 8'h00; 14'h03A2: rddata <= 8'h39; 14'h03A3: rddata <= 8'h7E;
            14'h03A4: rddata <= 8'h23; 14'h03A5: rddata <= 8'hFE; 14'h03A6: rddata <= 8'h81; 14'h03A7: rddata <= 8'hC0;
            14'h03A8: rddata <= 8'h4E; 14'h03A9: rddata <= 8'h23; 14'h03AA: rddata <= 8'h46; 14'h03AB: rddata <= 8'h23;
            14'h03AC: rddata <= 8'hE5; 14'h03AD: rddata <= 8'h60; 14'h03AE: rddata <= 8'h69; 14'h03AF: rddata <= 8'h7A;
            14'h03B0: rddata <= 8'hB3; 14'h03B1: rddata <= 8'hEB; 14'h03B2: rddata <= 8'h28; 14'h03B3: rddata <= 8'h02;
            14'h03B4: rddata <= 8'hEB; 14'h03B5: rddata <= 8'hE7; 14'h03B6: rddata <= 8'h01; 14'h03B7: rddata <= 8'h0D;
            14'h03B8: rddata <= 8'h00; 14'h03B9: rddata <= 8'hE1; 14'h03BA: rddata <= 8'hC8; 14'h03BB: rddata <= 8'h09;
            14'h03BC: rddata <= 8'h18; 14'h03BD: rddata <= 8'hE5; 14'h03BE: rddata <= 8'h2A; 14'h03BF: rddata <= 8'hC9;
            14'h03C0: rddata <= 8'h38; 14'h03C1: rddata <= 8'h22; 14'h03C2: rddata <= 8'h4D; 14'h03C3: rddata <= 8'h38;
            14'h03C4: rddata <= 8'h1E; 14'h03C5: rddata <= 8'h02; 14'h03C6: rddata <= 8'h01; 14'h03C7: rddata <= 8'h1E;
            14'h03C8: rddata <= 8'h14; 14'h03C9: rddata <= 8'h01; 14'h03CA: rddata <= 8'h1E; 14'h03CB: rddata <= 8'h00;
            14'h03CC: rddata <= 8'h01; 14'h03CD: rddata <= 8'h1E; 14'h03CE: rddata <= 8'h12; 14'h03CF: rddata <= 8'h01;
            14'h03D0: rddata <= 8'h1E; 14'h03D1: rddata <= 8'h22; 14'h03D2: rddata <= 8'h01; 14'h03D3: rddata <= 8'h1E;
            14'h03D4: rddata <= 8'h0A; 14'h03D5: rddata <= 8'h01; 14'h03D6: rddata <= 8'h1E; 14'h03D7: rddata <= 8'h24;
            14'h03D8: rddata <= 8'h01; 14'h03D9: rddata <= 8'h1E; 14'h03DA: rddata <= 8'h18; 14'h03DB: rddata <= 8'hCD;
            14'h03DC: rddata <= 8'hE5; 14'h03DD: rddata <= 8'h0B; 14'h03DE: rddata <= 8'hF7; 14'h03DF: rddata <= 8'h00;
            14'h03E0: rddata <= 8'hCD; 14'h03E1: rddata <= 8'hDE; 14'h03E2: rddata <= 8'h19; 14'h03E3: rddata <= 8'h21;
            14'h03E4: rddata <= 8'h79; 14'h03E5: rddata <= 8'h03; 14'h03E6: rddata <= 8'hF7; 14'h03E7: rddata <= 8'h01;
            14'h03E8: rddata <= 8'h57; 14'h03E9: rddata <= 8'h19; 14'h03EA: rddata <= 8'h3E; 14'h03EB: rddata <= 8'h3F;
            14'h03EC: rddata <= 8'hDF; 14'h03ED: rddata <= 8'h7E; 14'h03EE: rddata <= 8'hDF; 14'h03EF: rddata <= 8'hD7;
            14'h03F0: rddata <= 8'hDF; 14'h03F1: rddata <= 8'h21; 14'h03F2: rddata <= 8'h61; 14'h03F3: rddata <= 8'h03;
            14'h03F4: rddata <= 8'hCD; 14'h03F5: rddata <= 8'h9D; 14'h03F6: rddata <= 8'h0E; 14'h03F7: rddata <= 8'h2A;
            14'h03F8: rddata <= 8'h4D; 14'h03F9: rddata <= 8'h38; 14'h03FA: rddata <= 8'h7C; 14'h03FB: rddata <= 8'hA5;
            14'h03FC: rddata <= 8'h3C; 14'h03FD: rddata <= 8'hC4; 14'h03FE: rddata <= 8'h6D; 14'h03FF: rddata <= 8'h16;
            14'h0400: rddata <= 8'h3E; 14'h0401: rddata <= 8'hC1; 14'h0402: rddata <= 8'hF7; 14'h0403: rddata <= 8'h02;
            14'h0404: rddata <= 8'hCD; 14'h0405: rddata <= 8'hBE; 14'h0406: rddata <= 8'h19; 14'h0407: rddata <= 8'hAF;
            14'h0408: rddata <= 8'h32; 14'h0409: rddata <= 8'h08; 14'h040A: rddata <= 8'h38; 14'h040B: rddata <= 8'hCD;
            14'h040C: rddata <= 8'hDE; 14'h040D: rddata <= 8'h19; 14'h040E: rddata <= 8'h21; 14'h040F: rddata <= 8'h6E;
            14'h0410: rddata <= 8'h03; 14'h0411: rddata <= 8'hCD; 14'h0412: rddata <= 8'h9D; 14'h0413: rddata <= 8'h0E;
            14'h0414: rddata <= 8'h21; 14'h0415: rddata <= 8'hFF; 14'h0416: rddata <= 8'hFF; 14'h0417: rddata <= 8'h22;
            14'h0418: rddata <= 8'h4D; 14'h0419: rddata <= 8'h38; 14'h041A: rddata <= 8'hCD; 14'h041B: rddata <= 8'h85;
            14'h041C: rddata <= 8'h0D; 14'h041D: rddata <= 8'h38; 14'h041E: rddata <= 8'hF5; 14'h041F: rddata <= 8'hD7;
            14'h0420: rddata <= 8'h3C; 14'h0421: rddata <= 8'h3D; 14'h0422: rddata <= 8'h28; 14'h0423: rddata <= 8'hF0;
            14'h0424: rddata <= 8'hF5; 14'h0425: rddata <= 8'hCD; 14'h0426: rddata <= 8'h9C; 14'h0427: rddata <= 8'h06;
            14'h0428: rddata <= 8'hD5; 14'h0429: rddata <= 8'hCD; 14'h042A: rddata <= 8'hBC; 14'h042B: rddata <= 8'h04;
            14'h042C: rddata <= 8'h47; 14'h042D: rddata <= 8'hD1; 14'h042E: rddata <= 8'hF1; 14'h042F: rddata <= 8'hF7;
            14'h0430: rddata <= 8'h03; 14'h0431: rddata <= 8'hD2; 14'h0432: rddata <= 8'h4B; 14'h0433: rddata <= 8'h06;
            14'h0434: rddata <= 8'hD5; 14'h0435: rddata <= 8'hC5; 14'h0436: rddata <= 8'hAF; 14'h0437: rddata <= 8'h32;
            14'h0438: rddata <= 8'hCC; 14'h0439: rddata <= 8'h38; 14'h043A: rddata <= 8'hD7; 14'h043B: rddata <= 8'hB7;
            14'h043C: rddata <= 8'hF5; 14'h043D: rddata <= 8'hCD; 14'h043E: rddata <= 8'h9F; 14'h043F: rddata <= 8'h04;
            14'h0440: rddata <= 8'h38; 14'h0441: rddata <= 8'h06; 14'h0442: rddata <= 8'hF1; 14'h0443: rddata <= 8'hF5;
            14'h0444: rddata <= 8'hCA; 14'h0445: rddata <= 8'hF3; 14'h0446: rddata <= 8'h06; 14'h0447: rddata <= 8'hB7;
            14'h0448: rddata <= 8'hC5; 14'h0449: rddata <= 8'h30; 14'h044A: rddata <= 8'h10; 14'h044B: rddata <= 8'hEB;
            14'h044C: rddata <= 8'h2A; 14'h044D: rddata <= 8'hD6; 14'h044E: rddata <= 8'h38; 14'h044F: rddata <= 8'h1A;
            14'h0450: rddata <= 8'h02; 14'h0451: rddata <= 8'h03; 14'h0452: rddata <= 8'h13; 14'h0453: rddata <= 8'hE7;
            14'h0454: rddata <= 8'h20; 14'h0455: rddata <= 8'hF9; 14'h0456: rddata <= 8'h60; 14'h0457: rddata <= 8'h69;
            14'h0458: rddata <= 8'h22; 14'h0459: rddata <= 8'hD6; 14'h045A: rddata <= 8'h38; 14'h045B: rddata <= 8'hD1;
            14'h045C: rddata <= 8'hF1; 14'h045D: rddata <= 8'h28; 14'h045E: rddata <= 8'h21; 14'h045F: rddata <= 8'h2A;
            14'h0460: rddata <= 8'hD6; 14'h0461: rddata <= 8'h38; 14'h0462: rddata <= 8'hE3; 14'h0463: rddata <= 8'hC1;
            14'h0464: rddata <= 8'h09; 14'h0465: rddata <= 8'hE5; 14'h0466: rddata <= 8'hCD; 14'h0467: rddata <= 8'h92;
            14'h0468: rddata <= 8'h0B; 14'h0469: rddata <= 8'hE1; 14'h046A: rddata <= 8'h22; 14'h046B: rddata <= 8'hD6;
            14'h046C: rddata <= 8'h38; 14'h046D: rddata <= 8'hEB; 14'h046E: rddata <= 8'h74; 14'h046F: rddata <= 8'hD1;
            14'h0470: rddata <= 8'h23; 14'h0471: rddata <= 8'h23; 14'h0472: rddata <= 8'h73; 14'h0473: rddata <= 8'h23;
            14'h0474: rddata <= 8'h72; 14'h0475: rddata <= 8'h23; 14'h0476: rddata <= 8'h11; 14'h0477: rddata <= 8'h60;
            14'h0478: rddata <= 8'h38; 14'h0479: rddata <= 8'h1A; 14'h047A: rddata <= 8'h77; 14'h047B: rddata <= 8'h23;
            14'h047C: rddata <= 8'h13; 14'h047D: rddata <= 8'hB7; 14'h047E: rddata <= 8'h20; 14'h047F: rddata <= 8'hF9;
            14'h0480: rddata <= 8'hF7; 14'h0481: rddata <= 8'h04; 14'h0482: rddata <= 8'hCD; 14'h0483: rddata <= 8'hCB;
            14'h0484: rddata <= 8'h0B; 14'h0485: rddata <= 8'hF7; 14'h0486: rddata <= 8'h05; 14'h0487: rddata <= 8'h23;
            14'h0488: rddata <= 8'hEB; 14'h0489: rddata <= 8'h62; 14'h048A: rddata <= 8'h6B; 14'h048B: rddata <= 8'h7E;
            14'h048C: rddata <= 8'h23; 14'h048D: rddata <= 8'hB6; 14'h048E: rddata <= 8'hCA; 14'h048F: rddata <= 8'h14;
            14'h0490: rddata <= 8'h04; 14'h0491: rddata <= 8'h23; 14'h0492: rddata <= 8'h23; 14'h0493: rddata <= 8'h23;
            14'h0494: rddata <= 8'hAF; 14'h0495: rddata <= 8'hBE; 14'h0496: rddata <= 8'h23; 14'h0497: rddata <= 8'h20;
            14'h0498: rddata <= 8'hFC; 14'h0499: rddata <= 8'hEB; 14'h049A: rddata <= 8'h73; 14'h049B: rddata <= 8'h23;
            14'h049C: rddata <= 8'h72; 14'h049D: rddata <= 8'h18; 14'h049E: rddata <= 8'hEA; 14'h049F: rddata <= 8'h2A;
            14'h04A0: rddata <= 8'h4F; 14'h04A1: rddata <= 8'h38; 14'h04A2: rddata <= 8'h44; 14'h04A3: rddata <= 8'h4D;
            14'h04A4: rddata <= 8'h7E; 14'h04A5: rddata <= 8'h23; 14'h04A6: rddata <= 8'hB6; 14'h04A7: rddata <= 8'h2B;
            14'h04A8: rddata <= 8'hC8; 14'h04A9: rddata <= 8'h23; 14'h04AA: rddata <= 8'h23; 14'h04AB: rddata <= 8'h7E;
            14'h04AC: rddata <= 8'h23; 14'h04AD: rddata <= 8'h66; 14'h04AE: rddata <= 8'h6F; 14'h04AF: rddata <= 8'hE7;
            14'h04B0: rddata <= 8'h60; 14'h04B1: rddata <= 8'h69; 14'h04B2: rddata <= 8'h7E; 14'h04B3: rddata <= 8'h23;
            14'h04B4: rddata <= 8'h66; 14'h04B5: rddata <= 8'h6F; 14'h04B6: rddata <= 8'h3F; 14'h04B7: rddata <= 8'hC8;
            14'h04B8: rddata <= 8'h3F; 14'h04B9: rddata <= 8'hD0; 14'h04BA: rddata <= 8'h18; 14'h04BB: rddata <= 8'hE6;
            14'h04BC: rddata <= 8'hAF; 14'h04BD: rddata <= 8'h32; 14'h04BE: rddata <= 8'hAC; 14'h04BF: rddata <= 8'h38;
            14'h04C0: rddata <= 8'h0E; 14'h04C1: rddata <= 8'h05; 14'h04C2: rddata <= 8'h11; 14'h04C3: rddata <= 8'h60;
            14'h04C4: rddata <= 8'h38; 14'h04C5: rddata <= 8'h7E; 14'h04C6: rddata <= 8'hFE; 14'h04C7: rddata <= 8'h20;
            14'h04C8: rddata <= 8'hCA; 14'h04C9: rddata <= 8'h3C; 14'h04CA: rddata <= 8'h05; 14'h04CB: rddata <= 8'h47;
            14'h04CC: rddata <= 8'hFE; 14'h04CD: rddata <= 8'h22; 14'h04CE: rddata <= 8'hCA; 14'h04CF: rddata <= 8'h58;
            14'h04D0: rddata <= 8'h05; 14'h04D1: rddata <= 8'hB7; 14'h04D2: rddata <= 8'hCA; 14'h04D3: rddata <= 8'h5E;
            14'h04D4: rddata <= 8'h05; 14'h04D5: rddata <= 8'h3A; 14'h04D6: rddata <= 8'hAC; 14'h04D7: rddata <= 8'h38;
            14'h04D8: rddata <= 8'hB7; 14'h04D9: rddata <= 8'h7E; 14'h04DA: rddata <= 8'hC2; 14'h04DB: rddata <= 8'h3C;
            14'h04DC: rddata <= 8'h05; 14'h04DD: rddata <= 8'hFE; 14'h04DE: rddata <= 8'h3F; 14'h04DF: rddata <= 8'h3E;
            14'h04E0: rddata <= 8'h95; 14'h04E1: rddata <= 8'hCA; 14'h04E2: rddata <= 8'h3C; 14'h04E3: rddata <= 8'h05;
            14'h04E4: rddata <= 8'h7E; 14'h04E5: rddata <= 8'hFE; 14'h04E6: rddata <= 8'h30; 14'h04E7: rddata <= 8'h38;
            14'h04E8: rddata <= 8'h05; 14'h04E9: rddata <= 8'hFE; 14'h04EA: rddata <= 8'h3C; 14'h04EB: rddata <= 8'hDA;
            14'h04EC: rddata <= 8'h3C; 14'h04ED: rddata <= 8'h05; 14'h04EE: rddata <= 8'hD5; 14'h04EF: rddata <= 8'h11;
            14'h04F0: rddata <= 8'h44; 14'h04F1: rddata <= 8'h02; 14'h04F2: rddata <= 8'hC5; 14'h04F3: rddata <= 8'h01;
            14'h04F4: rddata <= 8'h36; 14'h04F5: rddata <= 8'h05; 14'h04F6: rddata <= 8'hC5; 14'h04F7: rddata <= 8'h06;
            14'h04F8: rddata <= 8'h7F; 14'h04F9: rddata <= 8'h7E; 14'h04FA: rddata <= 8'hFE; 14'h04FB: rddata <= 8'h61;
            14'h04FC: rddata <= 8'h38; 14'h04FD: rddata <= 8'h07; 14'h04FE: rddata <= 8'hFE; 14'h04FF: rddata <= 8'h7B;
            14'h0500: rddata <= 8'h30; 14'h0501: rddata <= 8'h03; 14'h0502: rddata <= 8'hE6; 14'h0503: rddata <= 8'h5F;
            14'h0504: rddata <= 8'h77; 14'h0505: rddata <= 8'h4E; 14'h0506: rddata <= 8'hEB; 14'h0507: rddata <= 8'h23;
            14'h0508: rddata <= 8'hB6; 14'h0509: rddata <= 8'hF2; 14'h050A: rddata <= 8'h07; 14'h050B: rddata <= 8'h05;
            14'h050C: rddata <= 8'h04; 14'h050D: rddata <= 8'h7E; 14'h050E: rddata <= 8'hE6; 14'h050F: rddata <= 8'h7F;
            14'h0510: rddata <= 8'hC8; 14'h0511: rddata <= 8'hB9; 14'h0512: rddata <= 8'h20; 14'h0513: rddata <= 8'hF3;
            14'h0514: rddata <= 8'hEB; 14'h0515: rddata <= 8'hE5; 14'h0516: rddata <= 8'h13; 14'h0517: rddata <= 8'h1A;
            14'h0518: rddata <= 8'hB7; 14'h0519: rddata <= 8'hFA; 14'h051A: rddata <= 8'h32; 14'h051B: rddata <= 8'h05;
            14'h051C: rddata <= 8'h4F; 14'h051D: rddata <= 8'h78; 14'h051E: rddata <= 8'hFE; 14'h051F: rddata <= 8'h88;
            14'h0520: rddata <= 8'h20; 14'h0521: rddata <= 8'h02; 14'h0522: rddata <= 8'hD7; 14'h0523: rddata <= 8'h2B;
            14'h0524: rddata <= 8'h23; 14'h0525: rddata <= 8'h7E; 14'h0526: rddata <= 8'hFE; 14'h0527: rddata <= 8'h61;
            14'h0528: rddata <= 8'h38; 14'h0529: rddata <= 8'h02; 14'h052A: rddata <= 8'hE6; 14'h052B: rddata <= 8'h5F;
            14'h052C: rddata <= 8'hB9; 14'h052D: rddata <= 8'h28; 14'h052E: rddata <= 8'hE7; 14'h052F: rddata <= 8'hE1;
            14'h0530: rddata <= 8'h18; 14'h0531: rddata <= 8'hD3; 14'h0532: rddata <= 8'h48; 14'h0533: rddata <= 8'hF1;
            14'h0534: rddata <= 8'hEB; 14'h0535: rddata <= 8'hC9; 14'h0536: rddata <= 8'hF7; 14'h0537: rddata <= 8'h0A;
            14'h0538: rddata <= 8'hEB; 14'h0539: rddata <= 8'h79; 14'h053A: rddata <= 8'hC1; 14'h053B: rddata <= 8'hD1;
            14'h053C: rddata <= 8'h23; 14'h053D: rddata <= 8'h12; 14'h053E: rddata <= 8'h13; 14'h053F: rddata <= 8'h0C;
            14'h0540: rddata <= 8'hD6; 14'h0541: rddata <= 8'h3A; 14'h0542: rddata <= 8'h28; 14'h0543: rddata <= 8'h04;
            14'h0544: rddata <= 8'hFE; 14'h0545: rddata <= 8'h49; 14'h0546: rddata <= 8'h20; 14'h0547: rddata <= 8'h03;
            14'h0548: rddata <= 8'h32; 14'h0549: rddata <= 8'hAC; 14'h054A: rddata <= 8'h38; 14'h054B: rddata <= 8'hD6;
            14'h054C: rddata <= 8'h54; 14'h054D: rddata <= 8'hC2; 14'h054E: rddata <= 8'hC5; 14'h054F: rddata <= 8'h04;
            14'h0550: rddata <= 8'h47; 14'h0551: rddata <= 8'h7E; 14'h0552: rddata <= 8'hB7; 14'h0553: rddata <= 8'h28;
            14'h0554: rddata <= 8'h09; 14'h0555: rddata <= 8'hB8; 14'h0556: rddata <= 8'h28; 14'h0557: rddata <= 8'hE4;
            14'h0558: rddata <= 8'h23; 14'h0559: rddata <= 8'h12; 14'h055A: rddata <= 8'h0C; 14'h055B: rddata <= 8'h13;
            14'h055C: rddata <= 8'h18; 14'h055D: rddata <= 8'hF3; 14'h055E: rddata <= 8'h21; 14'h055F: rddata <= 8'h5F;
            14'h0560: rddata <= 8'h38; 14'h0561: rddata <= 8'h12; 14'h0562: rddata <= 8'h13; 14'h0563: rddata <= 8'h12;
            14'h0564: rddata <= 8'h13; 14'h0565: rddata <= 8'h12; 14'h0566: rddata <= 8'hC9; 14'h0567: rddata <= 8'h3E;
            14'h0568: rddata <= 8'h01; 14'h0569: rddata <= 8'h32; 14'h056A: rddata <= 8'h47; 14'h056B: rddata <= 8'h38;
            14'h056C: rddata <= 8'h3E; 14'h056D: rddata <= 8'h17; 14'h056E: rddata <= 8'h32; 14'h056F: rddata <= 8'h08;
            14'h0570: rddata <= 8'h38; 14'h0571: rddata <= 8'hCD; 14'h0572: rddata <= 8'h9C; 14'h0573: rddata <= 8'h06;
            14'h0574: rddata <= 8'hC0; 14'h0575: rddata <= 8'hC1; 14'h0576: rddata <= 8'hCD; 14'h0577: rddata <= 8'h9F;
            14'h0578: rddata <= 8'h04; 14'h0579: rddata <= 8'hC5; 14'h057A: rddata <= 8'hE1; 14'h057B: rddata <= 8'h4E;
            14'h057C: rddata <= 8'h23; 14'h057D: rddata <= 8'h46; 14'h057E: rddata <= 8'h23; 14'h057F: rddata <= 8'h78;
            14'h0580: rddata <= 8'hB1; 14'h0581: rddata <= 8'hCA; 14'h0582: rddata <= 8'h02; 14'h0583: rddata <= 8'h04;
            14'h0584: rddata <= 8'hCD; 14'h0585: rddata <= 8'h25; 14'h0586: rddata <= 8'h1A; 14'h0587: rddata <= 8'hC5;
            14'h0588: rddata <= 8'hCD; 14'h0589: rddata <= 8'hEA; 14'h058A: rddata <= 8'h19; 14'h058B: rddata <= 8'h5E;
            14'h058C: rddata <= 8'h23; 14'h058D: rddata <= 8'h56; 14'h058E: rddata <= 8'h23; 14'h058F: rddata <= 8'hE5;
            14'h0590: rddata <= 8'hEB; 14'h0591: rddata <= 8'hCD; 14'h0592: rddata <= 8'h75; 14'h0593: rddata <= 8'h16;
            14'h0594: rddata <= 8'h3E; 14'h0595: rddata <= 8'h20; 14'h0596: rddata <= 8'hE1; 14'h0597: rddata <= 8'hDF;
            14'h0598: rddata <= 8'h7E; 14'h0599: rddata <= 8'h23; 14'h059A: rddata <= 8'hB7; 14'h059B: rddata <= 8'h28;
            14'h059C: rddata <= 8'hDD; 14'h059D: rddata <= 8'hF2; 14'h059E: rddata <= 8'h97; 14'h059F: rddata <= 8'h05;
            14'h05A0: rddata <= 8'hF7; 14'h05A1: rddata <= 8'h16; 14'h05A2: rddata <= 8'hD6; 14'h05A3: rddata <= 8'h7F;
            14'h05A4: rddata <= 8'h4F; 14'h05A5: rddata <= 8'h11; 14'h05A6: rddata <= 8'h45; 14'h05A7: rddata <= 8'h02;
            14'h05A8: rddata <= 8'h1A; 14'h05A9: rddata <= 8'h13; 14'h05AA: rddata <= 8'hB7; 14'h05AB: rddata <= 8'hF2;
            14'h05AC: rddata <= 8'hA8; 14'h05AD: rddata <= 8'h05; 14'h05AE: rddata <= 8'h0D; 14'h05AF: rddata <= 8'h20;
            14'h05B0: rddata <= 8'hF7; 14'h05B1: rddata <= 8'hE6; 14'h05B2: rddata <= 8'h7F; 14'h05B3: rddata <= 8'hDF;
            14'h05B4: rddata <= 8'h1A; 14'h05B5: rddata <= 8'h13; 14'h05B6: rddata <= 8'hB7; 14'h05B7: rddata <= 8'hF2;
            14'h05B8: rddata <= 8'hB1; 14'h05B9: rddata <= 8'h05; 14'h05BA: rddata <= 8'h18; 14'h05BB: rddata <= 8'hDC;
            14'h05BC: rddata <= 8'h3E; 14'h05BD: rddata <= 8'h64; 14'h05BE: rddata <= 8'h32; 14'h05BF: rddata <= 8'hCB;
            14'h05C0: rddata <= 8'h38; 14'h05C1: rddata <= 8'hCD; 14'h05C2: rddata <= 8'h31; 14'h05C3: rddata <= 8'h07;
            14'h05C4: rddata <= 8'hC1; 14'h05C5: rddata <= 8'hE5; 14'h05C6: rddata <= 8'hCD; 14'h05C7: rddata <= 8'h1C;
            14'h05C8: rddata <= 8'h07; 14'h05C9: rddata <= 8'h22; 14'h05CA: rddata <= 8'hC7; 14'h05CB: rddata <= 8'h38;
            14'h05CC: rddata <= 8'h21; 14'h05CD: rddata <= 8'h02; 14'h05CE: rddata <= 8'h00; 14'h05CF: rddata <= 8'h39;
            14'h05D0: rddata <= 8'hCD; 14'h05D1: rddata <= 8'hA3; 14'h05D2: rddata <= 8'h03; 14'h05D3: rddata <= 8'h20;
            14'h05D4: rddata <= 8'h14; 14'h05D5: rddata <= 8'h09; 14'h05D6: rddata <= 8'hD5; 14'h05D7: rddata <= 8'h2B;
            14'h05D8: rddata <= 8'h56; 14'h05D9: rddata <= 8'h2B; 14'h05DA: rddata <= 8'h5E; 14'h05DB: rddata <= 8'h23;
            14'h05DC: rddata <= 8'h23; 14'h05DD: rddata <= 8'hE5; 14'h05DE: rddata <= 8'h2A; 14'h05DF: rddata <= 8'hC7;
            14'h05E0: rddata <= 8'h38; 14'h05E1: rddata <= 8'hE7; 14'h05E2: rddata <= 8'hE1; 14'h05E3: rddata <= 8'hD1;
            14'h05E4: rddata <= 8'h20; 14'h05E5: rddata <= 8'hEA; 14'h05E6: rddata <= 8'hD1; 14'h05E7: rddata <= 8'hF9;
            14'h05E8: rddata <= 8'h0C; 14'h05E9: rddata <= 8'hD1; 14'h05EA: rddata <= 8'hEB; 14'h05EB: rddata <= 8'h0E;
            14'h05EC: rddata <= 8'h08; 14'h05ED: rddata <= 8'hCD; 14'h05EE: rddata <= 8'hA0; 14'h05EF: rddata <= 8'h0B;
            14'h05F0: rddata <= 8'hE5; 14'h05F1: rddata <= 8'h2A; 14'h05F2: rddata <= 8'hC7; 14'h05F3: rddata <= 8'h38;
            14'h05F4: rddata <= 8'hE3; 14'h05F5: rddata <= 8'hE5; 14'h05F6: rddata <= 8'h2A; 14'h05F7: rddata <= 8'h4D;
            14'h05F8: rddata <= 8'h38; 14'h05F9: rddata <= 8'hE3; 14'h05FA: rddata <= 8'hCD; 14'h05FB: rddata <= 8'h75;
            14'h05FC: rddata <= 8'h09; 14'h05FD: rddata <= 8'hCF; 14'h05FE: rddata <= 8'hA1; 14'h05FF: rddata <= 8'hCD;
            14'h0600: rddata <= 8'h72; 14'h0601: rddata <= 8'h09; 14'h0602: rddata <= 8'hE5; 14'h0603: rddata <= 8'hCD;
            14'h0604: rddata <= 8'h2E; 14'h0605: rddata <= 8'h15; 14'h0606: rddata <= 8'hE1; 14'h0607: rddata <= 8'hC5;
            14'h0608: rddata <= 8'hD5; 14'h0609: rddata <= 8'h01; 14'h060A: rddata <= 8'h00; 14'h060B: rddata <= 8'h81;
            14'h060C: rddata <= 8'h51; 14'h060D: rddata <= 8'h5A; 14'h060E: rddata <= 8'h7E; 14'h060F: rddata <= 8'hFE;
            14'h0610: rddata <= 8'hA7; 14'h0611: rddata <= 8'h3E; 14'h0612: rddata <= 8'h01; 14'h0613: rddata <= 8'h20;
            14'h0614: rddata <= 8'h0A; 14'h0615: rddata <= 8'hD7; 14'h0616: rddata <= 8'hCD; 14'h0617: rddata <= 8'h72;
            14'h0618: rddata <= 8'h09; 14'h0619: rddata <= 8'hE5; 14'h061A: rddata <= 8'hCD; 14'h061B: rddata <= 8'h2E;
            14'h061C: rddata <= 8'h15; 14'h061D: rddata <= 8'hEF; 14'h061E: rddata <= 8'hE1; 14'h061F: rddata <= 8'hC5;
            14'h0620: rddata <= 8'hD5; 14'h0621: rddata <= 8'hF5; 14'h0622: rddata <= 8'h33; 14'h0623: rddata <= 8'hE5;
            14'h0624: rddata <= 8'h2A; 14'h0625: rddata <= 8'hCE; 14'h0626: rddata <= 8'h38; 14'h0627: rddata <= 8'hE3;
            14'h0628: rddata <= 8'h06; 14'h0629: rddata <= 8'h81; 14'h062A: rddata <= 8'hC5; 14'h062B: rddata <= 8'h33;
            14'h062C: rddata <= 8'h22; 14'h062D: rddata <= 8'hCE; 14'h062E: rddata <= 8'h38; 14'h062F: rddata <= 8'hCD;
            14'h0630: rddata <= 8'hC2; 14'h0631: rddata <= 8'h1F; 14'h0632: rddata <= 8'h7E; 14'h0633: rddata <= 8'hFE;
            14'h0634: rddata <= 8'h3A; 14'h0635: rddata <= 8'h28; 14'h0636: rddata <= 8'h14; 14'h0637: rddata <= 8'hB7;
            14'h0638: rddata <= 8'hC2; 14'h0639: rddata <= 8'hC4; 14'h063A: rddata <= 8'h03; 14'h063B: rddata <= 8'h23;
            14'h063C: rddata <= 8'h7E; 14'h063D: rddata <= 8'h23; 14'h063E: rddata <= 8'hB6; 14'h063F: rddata <= 8'hCA;
            14'h0640: rddata <= 8'h29; 14'h0641: rddata <= 8'h0C; 14'h0642: rddata <= 8'h23; 14'h0643: rddata <= 8'h5E;
            14'h0644: rddata <= 8'h23; 14'h0645: rddata <= 8'h56; 14'h0646: rddata <= 8'hEB; 14'h0647: rddata <= 8'h22;
            14'h0648: rddata <= 8'h4D; 14'h0649: rddata <= 8'h38; 14'h064A: rddata <= 8'hEB; 14'h064B: rddata <= 8'hD7;
            14'h064C: rddata <= 8'h11; 14'h064D: rddata <= 8'h2C; 14'h064E: rddata <= 8'h06; 14'h064F: rddata <= 8'hD5;
            14'h0650: rddata <= 8'hC8; 14'h0651: rddata <= 8'hD6; 14'h0652: rddata <= 8'h80; 14'h0653: rddata <= 8'hDA;
            14'h0654: rddata <= 8'h31; 14'h0655: rddata <= 8'h07; 14'h0656: rddata <= 8'hFE; 14'h0657: rddata <= 8'h20;
            14'h0658: rddata <= 8'hF7; 14'h0659: rddata <= 8'h17; 14'h065A: rddata <= 8'hD2; 14'h065B: rddata <= 8'hC4;
            14'h065C: rddata <= 8'h03; 14'h065D: rddata <= 8'h07; 14'h065E: rddata <= 8'h4F; 14'h065F: rddata <= 8'h06;
            14'h0660: rddata <= 8'h00; 14'h0661: rddata <= 8'hEB; 14'h0662: rddata <= 8'h21; 14'h0663: rddata <= 8'hD5;
            14'h0664: rddata <= 8'h01; 14'h0665: rddata <= 8'h09; 14'h0666: rddata <= 8'h4E; 14'h0667: rddata <= 8'h23;
            14'h0668: rddata <= 8'h46; 14'h0669: rddata <= 8'hC5; 14'h066A: rddata <= 8'hEB; 14'h066B: rddata <= 8'h23;
            14'h066C: rddata <= 8'h7E; 14'h066D: rddata <= 8'hFE; 14'h066E: rddata <= 8'h3A; 14'h066F: rddata <= 8'hD0;
            14'h0670: rddata <= 8'hFE; 14'h0671: rddata <= 8'h20; 14'h0672: rddata <= 8'h28; 14'h0673: rddata <= 8'hF7;
            14'h0674: rddata <= 8'hFE; 14'h0675: rddata <= 8'h30; 14'h0676: rddata <= 8'h3F; 14'h0677: rddata <= 8'h3C;
            14'h0678: rddata <= 8'h3D; 14'h0679: rddata <= 8'hC9; 14'h067A: rddata <= 8'hD7; 14'h067B: rddata <= 8'hCD;
            14'h067C: rddata <= 8'h72; 14'h067D: rddata <= 8'h09; 14'h067E: rddata <= 8'hEF; 14'h067F: rddata <= 8'hFA;
            14'h0680: rddata <= 8'h97; 14'h0681: rddata <= 8'h06; 14'h0682: rddata <= 8'h3A; 14'h0683: rddata <= 8'hE7;
            14'h0684: rddata <= 8'h38; 14'h0685: rddata <= 8'hFE; 14'h0686: rddata <= 8'h90; 14'h0687: rddata <= 8'hDA;
            14'h0688: rddata <= 8'h86; 14'h0689: rddata <= 8'h15; 14'h068A: rddata <= 8'h01; 14'h068B: rddata <= 8'h80;
            14'h068C: rddata <= 8'h90; 14'h068D: rddata <= 8'h11; 14'h068E: rddata <= 8'h00; 14'h068F: rddata <= 8'h00;
            14'h0690: rddata <= 8'hE5; 14'h0691: rddata <= 8'hCD; 14'h0692: rddata <= 8'h5B; 14'h0693: rddata <= 8'h15;
            14'h0694: rddata <= 8'hE1; 14'h0695: rddata <= 8'h51; 14'h0696: rddata <= 8'hC8; 14'h0697: rddata <= 8'h1E;
            14'h0698: rddata <= 8'h08; 14'h0699: rddata <= 8'hC3; 14'h069A: rddata <= 8'hDB; 14'h069B: rddata <= 8'h03;
            14'h069C: rddata <= 8'h2B; 14'h069D: rddata <= 8'h11; 14'h069E: rddata <= 8'h00; 14'h069F: rddata <= 8'h00;
            14'h06A0: rddata <= 8'hD7; 14'h06A1: rddata <= 8'hD0; 14'h06A2: rddata <= 8'hE5; 14'h06A3: rddata <= 8'hF5;
            14'h06A4: rddata <= 8'h21; 14'h06A5: rddata <= 8'h98; 14'h06A6: rddata <= 8'h19; 14'h06A7: rddata <= 8'hE7;
            14'h06A8: rddata <= 8'h38; 14'h06A9: rddata <= 8'h11; 14'h06AA: rddata <= 8'h62; 14'h06AB: rddata <= 8'h6B;
            14'h06AC: rddata <= 8'h19; 14'h06AD: rddata <= 8'h29; 14'h06AE: rddata <= 8'h19; 14'h06AF: rddata <= 8'h29;
            14'h06B0: rddata <= 8'hF1; 14'h06B1: rddata <= 8'hD6; 14'h06B2: rddata <= 8'h30; 14'h06B3: rddata <= 8'h5F;
            14'h06B4: rddata <= 8'h16; 14'h06B5: rddata <= 8'h00; 14'h06B6: rddata <= 8'h19; 14'h06B7: rddata <= 8'hEB;
            14'h06B8: rddata <= 8'hE1; 14'h06B9: rddata <= 8'h18; 14'h06BA: rddata <= 8'hE5; 14'h06BB: rddata <= 8'hF1;
            14'h06BC: rddata <= 8'hE1; 14'h06BD: rddata <= 8'hC9; 14'h06BE: rddata <= 8'hF7; 14'h06BF: rddata <= 8'h18;
            14'h06C0: rddata <= 8'hCA; 14'h06C1: rddata <= 8'hCB; 14'h06C2: rddata <= 8'h0B; 14'h06C3: rddata <= 8'hCD;
            14'h06C4: rddata <= 8'hCF; 14'h06C5: rddata <= 8'h0B; 14'h06C6: rddata <= 8'h01; 14'h06C7: rddata <= 8'h2C;
            14'h06C8: rddata <= 8'h06; 14'h06C9: rddata <= 8'h18; 14'h06CA: rddata <= 8'h10; 14'h06CB: rddata <= 8'h0E;
            14'h06CC: rddata <= 8'h03; 14'h06CD: rddata <= 8'hCD; 14'h06CE: rddata <= 8'hA0; 14'h06CF: rddata <= 8'h0B;
            14'h06D0: rddata <= 8'hC1; 14'h06D1: rddata <= 8'hE5; 14'h06D2: rddata <= 8'hE5; 14'h06D3: rddata <= 8'h2A;
            14'h06D4: rddata <= 8'h4D; 14'h06D5: rddata <= 8'h38; 14'h06D6: rddata <= 8'hE3; 14'h06D7: rddata <= 8'h3E;
            14'h06D8: rddata <= 8'h8C; 14'h06D9: rddata <= 8'hF5; 14'h06DA: rddata <= 8'h33; 14'h06DB: rddata <= 8'hC5;
            14'h06DC: rddata <= 8'hCD; 14'h06DD: rddata <= 8'h9C; 14'h06DE: rddata <= 8'h06; 14'h06DF: rddata <= 8'hCD;
            14'h06E0: rddata <= 8'h1E; 14'h06E1: rddata <= 8'h07; 14'h06E2: rddata <= 8'h23; 14'h06E3: rddata <= 8'hE5;
            14'h06E4: rddata <= 8'h2A; 14'h06E5: rddata <= 8'h4D; 14'h06E6: rddata <= 8'h38; 14'h06E7: rddata <= 8'hE7;
            14'h06E8: rddata <= 8'hE1; 14'h06E9: rddata <= 8'hDC; 14'h06EA: rddata <= 8'hA2; 14'h06EB: rddata <= 8'h04;
            14'h06EC: rddata <= 8'hD4; 14'h06ED: rddata <= 8'h9F; 14'h06EE: rddata <= 8'h04; 14'h06EF: rddata <= 8'h60;
            14'h06F0: rddata <= 8'h69; 14'h06F1: rddata <= 8'h2B; 14'h06F2: rddata <= 8'hD8; 14'h06F3: rddata <= 8'h1E;
            14'h06F4: rddata <= 8'h0E; 14'h06F5: rddata <= 8'hC3; 14'h06F6: rddata <= 8'hDB; 14'h06F7: rddata <= 8'h03;
            14'h06F8: rddata <= 8'hC0; 14'h06F9: rddata <= 8'h16; 14'h06FA: rddata <= 8'hFF; 14'h06FB: rddata <= 8'hCD;
            14'h06FC: rddata <= 8'h9F; 14'h06FD: rddata <= 8'h03; 14'h06FE: rddata <= 8'hF9; 14'h06FF: rddata <= 8'hFE;
            14'h0700: rddata <= 8'h8C; 14'h0701: rddata <= 8'h1E; 14'h0702: rddata <= 8'h04; 14'h0703: rddata <= 8'hC2;
            14'h0704: rddata <= 8'hDB; 14'h0705: rddata <= 8'h03; 14'h0706: rddata <= 8'hE1; 14'h0707: rddata <= 8'h22;
            14'h0708: rddata <= 8'h4D; 14'h0709: rddata <= 8'h38; 14'h070A: rddata <= 8'h23; 14'h070B: rddata <= 8'h7C;
            14'h070C: rddata <= 8'hB5; 14'h070D: rddata <= 8'h20; 14'h070E: rddata <= 8'h07; 14'h070F: rddata <= 8'h3A;
            14'h0710: rddata <= 8'hCC; 14'h0711: rddata <= 8'h38; 14'h0712: rddata <= 8'hB7; 14'h0713: rddata <= 8'hC2;
            14'h0714: rddata <= 8'h01; 14'h0715: rddata <= 8'h04; 14'h0716: rddata <= 8'h21; 14'h0717: rddata <= 8'h2C;
            14'h0718: rddata <= 8'h06; 14'h0719: rddata <= 8'hE3; 14'h071A: rddata <= 8'h3E; 14'h071B: rddata <= 8'hE1;
            14'h071C: rddata <= 8'h01; 14'h071D: rddata <= 8'h3A; 14'h071E: rddata <= 8'h0E; 14'h071F: rddata <= 8'h00;
            14'h0720: rddata <= 8'h06; 14'h0721: rddata <= 8'h00; 14'h0722: rddata <= 8'h79; 14'h0723: rddata <= 8'h48;
            14'h0724: rddata <= 8'h47; 14'h0725: rddata <= 8'h7E; 14'h0726: rddata <= 8'hB7; 14'h0727: rddata <= 8'hC8;
            14'h0728: rddata <= 8'hB8; 14'h0729: rddata <= 8'hC8; 14'h072A: rddata <= 8'h23; 14'h072B: rddata <= 8'hFE;
            14'h072C: rddata <= 8'h22; 14'h072D: rddata <= 8'h28; 14'h072E: rddata <= 8'hF3; 14'h072F: rddata <= 8'h18;
            14'h0730: rddata <= 8'hF4; 14'h0731: rddata <= 8'hCD; 14'h0732: rddata <= 8'hD1; 14'h0733: rddata <= 8'h10;
            14'h0734: rddata <= 8'hCF; 14'h0735: rddata <= 8'hB0; 14'h0736: rddata <= 8'hD5; 14'h0737: rddata <= 8'h3A;
            14'h0738: rddata <= 8'hAB; 14'h0739: rddata <= 8'h38; 14'h073A: rddata <= 8'hF5; 14'h073B: rddata <= 8'hCD;
            14'h073C: rddata <= 8'h85; 14'h073D: rddata <= 8'h09; 14'h073E: rddata <= 8'hF1; 14'h073F: rddata <= 8'hE3;
            14'h0740: rddata <= 8'h22; 14'h0741: rddata <= 8'hCE; 14'h0742: rddata <= 8'h38; 14'h0743: rddata <= 8'h1F;
            14'h0744: rddata <= 8'hCD; 14'h0745: rddata <= 8'h77; 14'h0746: rddata <= 8'h09; 14'h0747: rddata <= 8'hCA;
            14'h0748: rddata <= 8'h79; 14'h0749: rddata <= 8'h07; 14'h074A: rddata <= 8'hE5; 14'h074B: rddata <= 8'h2A;
            14'h074C: rddata <= 8'hE4; 14'h074D: rddata <= 8'h38; 14'h074E: rddata <= 8'hE5; 14'h074F: rddata <= 8'h23;
            14'h0750: rddata <= 8'h23; 14'h0751: rddata <= 8'h5E; 14'h0752: rddata <= 8'h23; 14'h0753: rddata <= 8'h56;
            14'h0754: rddata <= 8'h2A; 14'h0755: rddata <= 8'h4F; 14'h0756: rddata <= 8'h38; 14'h0757: rddata <= 8'hE7;
            14'h0758: rddata <= 8'h30; 14'h0759: rddata <= 8'h0E; 14'h075A: rddata <= 8'h2A; 14'h075B: rddata <= 8'hDA;
            14'h075C: rddata <= 8'h38; 14'h075D: rddata <= 8'hE7; 14'h075E: rddata <= 8'hD1; 14'h075F: rddata <= 8'h30;
            14'h0760: rddata <= 8'h0F; 14'h0761: rddata <= 8'h21; 14'h0762: rddata <= 8'hBD; 14'h0763: rddata <= 8'h38;
            14'h0764: rddata <= 8'hE7; 14'h0765: rddata <= 8'h30; 14'h0766: rddata <= 8'h09; 14'h0767: rddata <= 8'h3E;
            14'h0768: rddata <= 8'hD1; 14'h0769: rddata <= 8'hCD; 14'h076A: rddata <= 8'hE4; 14'h076B: rddata <= 8'h0F;
            14'h076C: rddata <= 8'hEB; 14'h076D: rddata <= 8'hCD; 14'h076E: rddata <= 8'h39; 14'h076F: rddata <= 8'h0E;
            14'h0770: rddata <= 8'hCD; 14'h0771: rddata <= 8'hE4; 14'h0772: rddata <= 8'h0F; 14'h0773: rddata <= 8'hE1;
            14'h0774: rddata <= 8'hCD; 14'h0775: rddata <= 8'h3D; 14'h0776: rddata <= 8'h15; 14'h0777: rddata <= 8'hE1;
            14'h0778: rddata <= 8'hC9; 14'h0779: rddata <= 8'hE5; 14'h077A: rddata <= 8'hCD; 14'h077B: rddata <= 8'h3A;
            14'h077C: rddata <= 8'h15; 14'h077D: rddata <= 8'hD1; 14'h077E: rddata <= 8'hE1; 14'h077F: rddata <= 8'hC9;
            14'h0780: rddata <= 8'hF7; 14'h0781: rddata <= 8'h19; 14'h0782: rddata <= 8'hCD; 14'h0783: rddata <= 8'h54;
            14'h0784: rddata <= 8'h0B; 14'h0785: rddata <= 8'h7E; 14'h0786: rddata <= 8'h47; 14'h0787: rddata <= 8'hFE;
            14'h0788: rddata <= 8'h8C; 14'h0789: rddata <= 8'h28; 14'h078A: rddata <= 8'h03; 14'h078B: rddata <= 8'hCF;
            14'h078C: rddata <= 8'h88; 14'h078D: rddata <= 8'h2B; 14'h078E: rddata <= 8'h4B; 14'h078F: rddata <= 8'h0D;
            14'h0790: rddata <= 8'h78; 14'h0791: rddata <= 8'hCA; 14'h0792: rddata <= 8'h51; 14'h0793: rddata <= 8'h06;
            14'h0794: rddata <= 8'hCD; 14'h0795: rddata <= 8'h9D; 14'h0796: rddata <= 8'h06; 14'h0797: rddata <= 8'hFE;
            14'h0798: rddata <= 8'h2C; 14'h0799: rddata <= 8'hC0; 14'h079A: rddata <= 8'h18; 14'h079B: rddata <= 8'hF3;
            14'h079C: rddata <= 8'hCD; 14'h079D: rddata <= 8'h85; 14'h079E: rddata <= 8'h09; 14'h079F: rddata <= 8'h7E;
            14'h07A0: rddata <= 8'hFE; 14'h07A1: rddata <= 8'h88; 14'h07A2: rddata <= 8'h28; 14'h07A3: rddata <= 8'h03;
            14'h07A4: rddata <= 8'hCF; 14'h07A5: rddata <= 8'hA5; 14'h07A6: rddata <= 8'h2B; 14'h07A7: rddata <= 8'hCD;
            14'h07A8: rddata <= 8'h75; 14'h07A9: rddata <= 8'h09; 14'h07AA: rddata <= 8'hEF; 14'h07AB: rddata <= 8'hCA;
            14'h07AC: rddata <= 8'h1E; 14'h07AD: rddata <= 8'h07; 14'h07AE: rddata <= 8'hD7; 14'h07AF: rddata <= 8'hDA;
            14'h07B0: rddata <= 8'hDC; 14'h07B1: rddata <= 8'h06; 14'h07B2: rddata <= 8'hC3; 14'h07B3: rddata <= 8'h50;
            14'h07B4: rddata <= 8'h06; 14'h07B5: rddata <= 8'h3E; 14'h07B6: rddata <= 8'h01; 14'h07B7: rddata <= 8'h32;
            14'h07B8: rddata <= 8'h47; 14'h07B9: rddata <= 8'h38; 14'h07BA: rddata <= 8'h2B; 14'h07BB: rddata <= 8'hD7;
            14'h07BC: rddata <= 8'hF7; 14'h07BD: rddata <= 8'h06; 14'h07BE: rddata <= 8'hCC; 14'h07BF: rddata <= 8'hEA;
            14'h07C0: rddata <= 8'h19; 14'h07C1: rddata <= 8'hCA; 14'h07C2: rddata <= 8'h66; 14'h07C3: rddata <= 8'h08;
            14'h07C4: rddata <= 8'hFE; 14'h07C5: rddata <= 8'hA0; 14'h07C6: rddata <= 8'hCA; 14'h07C7: rddata <= 8'h3A;
            14'h07C8: rddata <= 8'h08; 14'h07C9: rddata <= 8'hFE; 14'h07CA: rddata <= 8'hA3; 14'h07CB: rddata <= 8'hCA;
            14'h07CC: rddata <= 8'h3A; 14'h07CD: rddata <= 8'h08; 14'h07CE: rddata <= 8'hE5; 14'h07CF: rddata <= 8'hFE;
            14'h07D0: rddata <= 8'h2C; 14'h07D1: rddata <= 8'h28; 14'h07D2: rddata <= 8'h44; 14'h07D3: rddata <= 8'hFE;
            14'h07D4: rddata <= 8'h3B; 14'h07D5: rddata <= 8'hCA; 14'h07D6: rddata <= 8'h61; 14'h07D7: rddata <= 8'h08;
            14'h07D8: rddata <= 8'hC1; 14'h07D9: rddata <= 8'hCD; 14'h07DA: rddata <= 8'h85; 14'h07DB: rddata <= 8'h09;
            14'h07DC: rddata <= 8'hE5; 14'h07DD: rddata <= 8'h3A; 14'h07DE: rddata <= 8'hAB; 14'h07DF: rddata <= 8'h38;
            14'h07E0: rddata <= 8'hB7; 14'h07E1: rddata <= 8'hC2; 14'h07E2: rddata <= 8'h11; 14'h07E3: rddata <= 8'h08;
            14'h07E4: rddata <= 8'hCD; 14'h07E5: rddata <= 8'h80; 14'h07E6: rddata <= 8'h16; 14'h07E7: rddata <= 8'hCD;
            14'h07E8: rddata <= 8'h5F; 14'h07E9: rddata <= 8'h0E; 14'h07EA: rddata <= 8'h36; 14'h07EB: rddata <= 8'h20;
            14'h07EC: rddata <= 8'h2A; 14'h07ED: rddata <= 8'hE4; 14'h07EE: rddata <= 8'h38; 14'h07EF: rddata <= 8'h3A;
            14'h07F0: rddata <= 8'h47; 14'h07F1: rddata <= 8'h38; 14'h07F2: rddata <= 8'hB7; 14'h07F3: rddata <= 8'h28;
            14'h07F4: rddata <= 8'h08; 14'h07F5: rddata <= 8'h3A; 14'h07F6: rddata <= 8'h46; 14'h07F7: rddata <= 8'h38;
            14'h07F8: rddata <= 8'h86; 14'h07F9: rddata <= 8'hFE; 14'h07FA: rddata <= 8'h84; 14'h07FB: rddata <= 8'h18;
            14'h07FC: rddata <= 8'h0D; 14'h07FD: rddata <= 8'h3A; 14'h07FE: rddata <= 8'h48; 14'h07FF: rddata <= 8'h38;
            14'h0800: rddata <= 8'h47; 14'h0801: rddata <= 8'h3C; 14'h0802: rddata <= 8'h28; 14'h0803: rddata <= 8'h09;
            14'h0804: rddata <= 8'h3A; 14'h0805: rddata <= 8'h00; 14'h0806: rddata <= 8'h38; 14'h0807: rddata <= 8'h86;
            14'h0808: rddata <= 8'h3D; 14'h0809: rddata <= 8'hB8; 14'h080A: rddata <= 8'hD4; 14'h080B: rddata <= 8'hEA;
            14'h080C: rddata <= 8'h19; 14'h080D: rddata <= 8'hCD; 14'h080E: rddata <= 8'hA0; 14'h080F: rddata <= 8'h0E;
            14'h0810: rddata <= 8'hAF; 14'h0811: rddata <= 8'hC4; 14'h0812: rddata <= 8'hA0; 14'h0813: rddata <= 8'h0E;
            14'h0814: rddata <= 8'hE1; 14'h0815: rddata <= 8'h18; 14'h0816: rddata <= 8'hA3; 14'h0817: rddata <= 8'h3A;
            14'h0818: rddata <= 8'h47; 14'h0819: rddata <= 8'h38; 14'h081A: rddata <= 8'hB7; 14'h081B: rddata <= 8'h28;
            14'h081C: rddata <= 8'h08; 14'h081D: rddata <= 8'h3A; 14'h081E: rddata <= 8'h46; 14'h081F: rddata <= 8'h38;
            14'h0820: rddata <= 8'hFE; 14'h0821: rddata <= 8'h70; 14'h0822: rddata <= 8'hC3; 14'h0823: rddata <= 8'h2D;
            14'h0824: rddata <= 8'h08; 14'h0825: rddata <= 8'h3A; 14'h0826: rddata <= 8'h49; 14'h0827: rddata <= 8'h38;
            14'h0828: rddata <= 8'h47; 14'h0829: rddata <= 8'h3A; 14'h082A: rddata <= 8'h00; 14'h082B: rddata <= 8'h38;
            14'h082C: rddata <= 8'hB8; 14'h082D: rddata <= 8'hD4; 14'h082E: rddata <= 8'hEA; 14'h082F: rddata <= 8'h19;
            14'h0830: rddata <= 8'hD2; 14'h0831: rddata <= 8'h61; 14'h0832: rddata <= 8'h08; 14'h0833: rddata <= 8'hD6;
            14'h0834: rddata <= 8'h0E; 14'h0835: rddata <= 8'h30; 14'h0836: rddata <= 8'hFC; 14'h0837: rddata <= 8'h2F;
            14'h0838: rddata <= 8'h18; 14'h0839: rddata <= 8'h20; 14'h083A: rddata <= 8'hF5; 14'h083B: rddata <= 8'hCD;
            14'h083C: rddata <= 8'h53; 14'h083D: rddata <= 8'h0B; 14'h083E: rddata <= 8'hCF; 14'h083F: rddata <= 8'h29;
            14'h0840: rddata <= 8'h2B; 14'h0841: rddata <= 8'hF1; 14'h0842: rddata <= 8'hD6; 14'h0843: rddata <= 8'hA3;
            14'h0844: rddata <= 8'hE5; 14'h0845: rddata <= 8'h28; 14'h0846: rddata <= 8'h0F; 14'h0847: rddata <= 8'h3A;
            14'h0848: rddata <= 8'h47; 14'h0849: rddata <= 8'h38; 14'h084A: rddata <= 8'hB7; 14'h084B: rddata <= 8'hCA;
            14'h084C: rddata <= 8'h53; 14'h084D: rddata <= 8'h08; 14'h084E: rddata <= 8'h3A; 14'h084F: rddata <= 8'h46;
            14'h0850: rddata <= 8'h38; 14'h0851: rddata <= 8'h18; 14'h0852: rddata <= 8'h03; 14'h0853: rddata <= 8'h3A;
            14'h0854: rddata <= 8'h00; 14'h0855: rddata <= 8'h38; 14'h0856: rddata <= 8'h2F; 14'h0857: rddata <= 8'h83;
            14'h0858: rddata <= 8'h30; 14'h0859: rddata <= 8'h07; 14'h085A: rddata <= 8'h3C; 14'h085B: rddata <= 8'h47;
            14'h085C: rddata <= 8'h3E; 14'h085D: rddata <= 8'h20; 14'h085E: rddata <= 8'hDF; 14'h085F: rddata <= 8'h10;
            14'h0860: rddata <= 8'hFD; 14'h0861: rddata <= 8'hE1; 14'h0862: rddata <= 8'hD7; 14'h0863: rddata <= 8'hC3;
            14'h0864: rddata <= 8'hC1; 14'h0865: rddata <= 8'h07; 14'h0866: rddata <= 8'hF7; 14'h0867: rddata <= 8'h07;
            14'h0868: rddata <= 8'hAF; 14'h0869: rddata <= 8'h32; 14'h086A: rddata <= 8'h47; 14'h086B: rddata <= 8'h38;
            14'h086C: rddata <= 8'hC9; 14'h086D: rddata <= 8'h3F; 14'h086E: rddata <= 8'h52; 14'h086F: rddata <= 8'h65;
            14'h0870: rddata <= 8'h64; 14'h0871: rddata <= 8'h6F; 14'h0872: rddata <= 8'h20; 14'h0873: rddata <= 8'h66;
            14'h0874: rddata <= 8'h72; 14'h0875: rddata <= 8'h6F; 14'h0876: rddata <= 8'h6D; 14'h0877: rddata <= 8'h20;
            14'h0878: rddata <= 8'h73; 14'h0879: rddata <= 8'h74; 14'h087A: rddata <= 8'h61; 14'h087B: rddata <= 8'h72;
            14'h087C: rddata <= 8'h74; 14'h087D: rddata <= 8'h0D; 14'h087E: rddata <= 8'h0A; 14'h087F: rddata <= 8'h00;
            14'h0880: rddata <= 8'hF7; 14'h0881: rddata <= 8'h08; 14'h0882: rddata <= 8'h3A; 14'h0883: rddata <= 8'hCD;
            14'h0884: rddata <= 8'h38; 14'h0885: rddata <= 8'hB7; 14'h0886: rddata <= 8'hC2; 14'h0887: rddata <= 8'hBE;
            14'h0888: rddata <= 8'h03; 14'h0889: rddata <= 8'hC1; 14'h088A: rddata <= 8'h21; 14'h088B: rddata <= 8'h6D;
            14'h088C: rddata <= 8'h08; 14'h088D: rddata <= 8'hCD; 14'h088E: rddata <= 8'h9D; 14'h088F: rddata <= 8'h0E;
            14'h0890: rddata <= 8'hC3; 14'h0891: rddata <= 8'h01; 14'h0892: rddata <= 8'h0C; 14'h0893: rddata <= 8'hF7;
            14'h0894: rddata <= 8'h1A; 14'h0895: rddata <= 8'hCD; 14'h0896: rddata <= 8'h45; 14'h0897: rddata <= 8'h0B;
            14'h0898: rddata <= 8'h7E; 14'h0899: rddata <= 8'hFE; 14'h089A: rddata <= 8'h22; 14'h089B: rddata <= 8'h3E;
            14'h089C: rddata <= 8'h00; 14'h089D: rddata <= 8'hC2; 14'h089E: rddata <= 8'hAA; 14'h089F: rddata <= 8'h08;
            14'h08A0: rddata <= 8'hCD; 14'h08A1: rddata <= 8'h60; 14'h08A2: rddata <= 8'h0E; 14'h08A3: rddata <= 8'hCF;
            14'h08A4: rddata <= 8'h3B; 14'h08A5: rddata <= 8'hE5; 14'h08A6: rddata <= 8'hCD; 14'h08A7: rddata <= 8'hA0;
            14'h08A8: rddata <= 8'h0E; 14'h08A9: rddata <= 8'h3E; 14'h08AA: rddata <= 8'hE5; 14'h08AB: rddata <= 8'hCD;
            14'h08AC: rddata <= 8'h5B; 14'h08AD: rddata <= 8'h0D; 14'h08AE: rddata <= 8'hC1; 14'h08AF: rddata <= 8'hDA;
            14'h08B0: rddata <= 8'h26; 14'h08B1: rddata <= 8'h0C; 14'h08B2: rddata <= 8'h23; 14'h08B3: rddata <= 8'h7E;
            14'h08B4: rddata <= 8'hB7; 14'h08B5: rddata <= 8'h2B; 14'h08B6: rddata <= 8'hC5; 14'h08B7: rddata <= 8'hCA;
            14'h08B8: rddata <= 8'h1B; 14'h08B9: rddata <= 8'h07; 14'h08BA: rddata <= 8'h36; 14'h08BB: rddata <= 8'h2C;
            14'h08BC: rddata <= 8'h18; 14'h08BD: rddata <= 8'h05; 14'h08BE: rddata <= 8'hE5; 14'h08BF: rddata <= 8'h2A;
            14'h08C0: rddata <= 8'hDC; 14'h08C1: rddata <= 8'h38; 14'h08C2: rddata <= 8'hF6; 14'h08C3: rddata <= 8'hAF;
            14'h08C4: rddata <= 8'h32; 14'h08C5: rddata <= 8'hCD; 14'h08C6: rddata <= 8'h38; 14'h08C7: rddata <= 8'hE3;
            14'h08C8: rddata <= 8'h01; 14'h08C9: rddata <= 8'hCF; 14'h08CA: rddata <= 8'h2C; 14'h08CB: rddata <= 8'hCD;
            14'h08CC: rddata <= 8'hD1; 14'h08CD: rddata <= 8'h10; 14'h08CE: rddata <= 8'hE3; 14'h08CF: rddata <= 8'hD5;
            14'h08D0: rddata <= 8'h7E; 14'h08D1: rddata <= 8'hFE; 14'h08D2: rddata <= 8'h2C; 14'h08D3: rddata <= 8'h28;
            14'h08D4: rddata <= 8'h1B; 14'h08D5: rddata <= 8'h3A; 14'h08D6: rddata <= 8'hCD; 14'h08D7: rddata <= 8'h38;
            14'h08D8: rddata <= 8'hB7; 14'h08D9: rddata <= 8'hC2; 14'h08DA: rddata <= 8'h53; 14'h08DB: rddata <= 8'h09;
            14'h08DC: rddata <= 8'h3E; 14'h08DD: rddata <= 8'h3F; 14'h08DE: rddata <= 8'hDF; 14'h08DF: rddata <= 8'hCD;
            14'h08E0: rddata <= 8'h5B; 14'h08E1: rddata <= 8'h0D; 14'h08E2: rddata <= 8'hD1; 14'h08E3: rddata <= 8'hC1;
            14'h08E4: rddata <= 8'hDA; 14'h08E5: rddata <= 8'h26; 14'h08E6: rddata <= 8'h0C; 14'h08E7: rddata <= 8'h23;
            14'h08E8: rddata <= 8'h7E; 14'h08E9: rddata <= 8'h2B; 14'h08EA: rddata <= 8'hB7; 14'h08EB: rddata <= 8'hC5;
            14'h08EC: rddata <= 8'hCA; 14'h08ED: rddata <= 8'h1B; 14'h08EE: rddata <= 8'h07; 14'h08EF: rddata <= 8'hD5;
            14'h08F0: rddata <= 8'hF7; 14'h08F1: rddata <= 8'h1C; 14'h08F2: rddata <= 8'h3A; 14'h08F3: rddata <= 8'hAB;
            14'h08F4: rddata <= 8'h38; 14'h08F5: rddata <= 8'hB7; 14'h08F6: rddata <= 8'h28; 14'h08F7: rddata <= 8'h1F;
            14'h08F8: rddata <= 8'hD7; 14'h08F9: rddata <= 8'h57; 14'h08FA: rddata <= 8'h47; 14'h08FB: rddata <= 8'hFE;
            14'h08FC: rddata <= 8'h22; 14'h08FD: rddata <= 8'h28; 14'h08FE: rddata <= 8'h0C; 14'h08FF: rddata <= 8'h3A;
            14'h0900: rddata <= 8'hCD; 14'h0901: rddata <= 8'h38; 14'h0902: rddata <= 8'hB7; 14'h0903: rddata <= 8'h57;
            14'h0904: rddata <= 8'h28; 14'h0905: rddata <= 8'h02; 14'h0906: rddata <= 8'h16; 14'h0907: rddata <= 8'h3A;
            14'h0908: rddata <= 8'h06; 14'h0909: rddata <= 8'h2C; 14'h090A: rddata <= 8'h2B; 14'h090B: rddata <= 8'hCD;
            14'h090C: rddata <= 8'h63; 14'h090D: rddata <= 8'h0E; 14'h090E: rddata <= 8'hEB; 14'h090F: rddata <= 8'h21;
            14'h0910: rddata <= 8'h20; 14'h0911: rddata <= 8'h09; 14'h0912: rddata <= 8'hE3; 14'h0913: rddata <= 8'hD5;
            14'h0914: rddata <= 8'hC3; 14'h0915: rddata <= 8'h4A; 14'h0916: rddata <= 8'h07; 14'h0917: rddata <= 8'hD7;
            14'h0918: rddata <= 8'hCD; 14'h0919: rddata <= 8'hE5; 14'h091A: rddata <= 8'h15; 14'h091B: rddata <= 8'hE3;
            14'h091C: rddata <= 8'hCD; 14'h091D: rddata <= 8'h3A; 14'h091E: rddata <= 8'h15; 14'h091F: rddata <= 8'hE1;
            14'h0920: rddata <= 8'h2B; 14'h0921: rddata <= 8'hD7; 14'h0922: rddata <= 8'h28; 14'h0923: rddata <= 8'h05;
            14'h0924: rddata <= 8'hFE; 14'h0925: rddata <= 8'h2C; 14'h0926: rddata <= 8'hC2; 14'h0927: rddata <= 8'h80;
            14'h0928: rddata <= 8'h08; 14'h0929: rddata <= 8'hE3; 14'h092A: rddata <= 8'h2B; 14'h092B: rddata <= 8'hD7;
            14'h092C: rddata <= 8'hC2; 14'h092D: rddata <= 8'hC9; 14'h092E: rddata <= 8'h08; 14'h092F: rddata <= 8'hD1;
            14'h0930: rddata <= 8'h3A; 14'h0931: rddata <= 8'hCD; 14'h0932: rddata <= 8'h38; 14'h0933: rddata <= 8'hB7;
            14'h0934: rddata <= 8'hEB; 14'h0935: rddata <= 8'hC2; 14'h0936: rddata <= 8'h1A; 14'h0937: rddata <= 8'h0C;
            14'h0938: rddata <= 8'hD5; 14'h0939: rddata <= 8'hB6; 14'h093A: rddata <= 8'h21; 14'h093B: rddata <= 8'h42;
            14'h093C: rddata <= 8'h09; 14'h093D: rddata <= 8'hC4; 14'h093E: rddata <= 8'h9D; 14'h093F: rddata <= 8'h0E;
            14'h0940: rddata <= 8'hE1; 14'h0941: rddata <= 8'hC9; 14'h0942: rddata <= 8'h3F; 14'h0943: rddata <= 8'h45;
            14'h0944: rddata <= 8'h78; 14'h0945: rddata <= 8'h74; 14'h0946: rddata <= 8'h72; 14'h0947: rddata <= 8'h61;
            14'h0948: rddata <= 8'h20; 14'h0949: rddata <= 8'h69; 14'h094A: rddata <= 8'h67; 14'h094B: rddata <= 8'h6E;
            14'h094C: rddata <= 8'h6F; 14'h094D: rddata <= 8'h72; 14'h094E: rddata <= 8'h65; 14'h094F: rddata <= 8'h64;
            14'h0950: rddata <= 8'h0D; 14'h0951: rddata <= 8'h0A; 14'h0952: rddata <= 8'h00; 14'h0953: rddata <= 8'hCD;
            14'h0954: rddata <= 8'h1C; 14'h0955: rddata <= 8'h07; 14'h0956: rddata <= 8'hB7; 14'h0957: rddata <= 8'h20;
            14'h0958: rddata <= 8'h11; 14'h0959: rddata <= 8'h23; 14'h095A: rddata <= 8'h7E; 14'h095B: rddata <= 8'h23;
            14'h095C: rddata <= 8'hB6; 14'h095D: rddata <= 8'h1E; 14'h095E: rddata <= 8'h06; 14'h095F: rddata <= 8'hCA;
            14'h0960: rddata <= 8'hDB; 14'h0961: rddata <= 8'h03; 14'h0962: rddata <= 8'h23; 14'h0963: rddata <= 8'h5E;
            14'h0964: rddata <= 8'h23; 14'h0965: rddata <= 8'h56; 14'h0966: rddata <= 8'hED; 14'h0967: rddata <= 8'h53;
            14'h0968: rddata <= 8'hC9; 14'h0969: rddata <= 8'h38; 14'h096A: rddata <= 8'hD7; 14'h096B: rddata <= 8'hFE;
            14'h096C: rddata <= 8'h83; 14'h096D: rddata <= 8'h20; 14'h096E: rddata <= 8'hE4; 14'h096F: rddata <= 8'hC3;
            14'h0970: rddata <= 8'hF0; 14'h0971: rddata <= 8'h08; 14'h0972: rddata <= 8'hCD; 14'h0973: rddata <= 8'h85;
            14'h0974: rddata <= 8'h09; 14'h0975: rddata <= 8'hF6; 14'h0976: rddata <= 8'h37; 14'h0977: rddata <= 8'h3A;
            14'h0978: rddata <= 8'hAB; 14'h0979: rddata <= 8'h38; 14'h097A: rddata <= 8'h8F; 14'h097B: rddata <= 8'hB7;
            14'h097C: rddata <= 8'hE8; 14'h097D: rddata <= 8'hC3; 14'h097E: rddata <= 8'hD9; 14'h097F: rddata <= 8'h03;
            14'h0980: rddata <= 8'hCF; 14'h0981: rddata <= 8'hB0; 14'h0982: rddata <= 8'h01; 14'h0983: rddata <= 8'hCF;
            14'h0984: rddata <= 8'h28; 14'h0985: rddata <= 8'h2B; 14'h0986: rddata <= 8'h16; 14'h0987: rddata <= 8'h00;
            14'h0988: rddata <= 8'hD5; 14'h0989: rddata <= 8'h0E; 14'h098A: rddata <= 8'h01; 14'h098B: rddata <= 8'hCD;
            14'h098C: rddata <= 8'hA0; 14'h098D: rddata <= 8'h0B; 14'h098E: rddata <= 8'hCD; 14'h098F: rddata <= 8'hFD;
            14'h0990: rddata <= 8'h09; 14'h0991: rddata <= 8'h22; 14'h0992: rddata <= 8'hD0; 14'h0993: rddata <= 8'h38;
            14'h0994: rddata <= 8'h2A; 14'h0995: rddata <= 8'hD0; 14'h0996: rddata <= 8'h38; 14'h0997: rddata <= 8'hC1;
            14'h0998: rddata <= 8'h78; 14'h0999: rddata <= 8'hFE; 14'h099A: rddata <= 8'h78; 14'h099B: rddata <= 8'hD4;
            14'h099C: rddata <= 8'h75; 14'h099D: rddata <= 8'h09; 14'h099E: rddata <= 8'h7E; 14'h099F: rddata <= 8'h22;
            14'h09A0: rddata <= 8'hC3; 14'h09A1: rddata <= 8'h38; 14'h09A2: rddata <= 8'hFE; 14'h09A3: rddata <= 8'hA8;
            14'h09A4: rddata <= 8'hD8; 14'h09A5: rddata <= 8'hFE; 14'h09A6: rddata <= 8'hB2; 14'h09A7: rddata <= 8'hD0;
            14'h09A8: rddata <= 8'hFE; 14'h09A9: rddata <= 8'hAF; 14'h09AA: rddata <= 8'hD2; 14'h09AB: rddata <= 8'hE2;
            14'h09AC: rddata <= 8'h09; 14'h09AD: rddata <= 8'hD6; 14'h09AE: rddata <= 8'hA8; 14'h09AF: rddata <= 8'h5F;
            14'h09B0: rddata <= 8'h20; 14'h09B1: rddata <= 8'h08; 14'h09B2: rddata <= 8'h3A; 14'h09B3: rddata <= 8'hAB;
            14'h09B4: rddata <= 8'h38; 14'h09B5: rddata <= 8'h3D; 14'h09B6: rddata <= 8'h7B; 14'h09B7: rddata <= 8'hCA;
            14'h09B8: rddata <= 8'h7C; 14'h09B9: rddata <= 8'h0F; 14'h09BA: rddata <= 8'h07; 14'h09BB: rddata <= 8'h83;
            14'h09BC: rddata <= 8'h5F; 14'h09BD: rddata <= 8'h21; 14'h09BE: rddata <= 8'h4C; 14'h09BF: rddata <= 8'h03;
            14'h09C0: rddata <= 8'h16; 14'h09C1: rddata <= 8'h00; 14'h09C2: rddata <= 8'h19; 14'h09C3: rddata <= 8'h78;
            14'h09C4: rddata <= 8'h56; 14'h09C5: rddata <= 8'hBA; 14'h09C6: rddata <= 8'hD0; 14'h09C7: rddata <= 8'h23;
            14'h09C8: rddata <= 8'hCD; 14'h09C9: rddata <= 8'h75; 14'h09CA: rddata <= 8'h09; 14'h09CB: rddata <= 8'hC5;
            14'h09CC: rddata <= 8'h01; 14'h09CD: rddata <= 8'h94; 14'h09CE: rddata <= 8'h09; 14'h09CF: rddata <= 8'hC5;
            14'h09D0: rddata <= 8'h43; 14'h09D1: rddata <= 8'h4A; 14'h09D2: rddata <= 8'hCD; 14'h09D3: rddata <= 8'h13;
            14'h09D4: rddata <= 8'h15; 14'h09D5: rddata <= 8'h58; 14'h09D6: rddata <= 8'h51; 14'h09D7: rddata <= 8'h4E;
            14'h09D8: rddata <= 8'h23; 14'h09D9: rddata <= 8'h46; 14'h09DA: rddata <= 8'h23; 14'h09DB: rddata <= 8'hC5;
            14'h09DC: rddata <= 8'h2A; 14'h09DD: rddata <= 8'hC3; 14'h09DE: rddata <= 8'h38; 14'h09DF: rddata <= 8'hC3;
            14'h09E0: rddata <= 8'h88; 14'h09E1: rddata <= 8'h09; 14'h09E2: rddata <= 8'h16; 14'h09E3: rddata <= 8'h00;
            14'h09E4: rddata <= 8'hD6; 14'h09E5: rddata <= 8'hAF; 14'h09E6: rddata <= 8'hDA; 14'h09E7: rddata <= 8'hD0;
            14'h09E8: rddata <= 8'h0A; 14'h09E9: rddata <= 8'hFE; 14'h09EA: rddata <= 8'h03; 14'h09EB: rddata <= 8'hD2;
            14'h09EC: rddata <= 8'hD0; 14'h09ED: rddata <= 8'h0A; 14'h09EE: rddata <= 8'hFE; 14'h09EF: rddata <= 8'h01;
            14'h09F0: rddata <= 8'h17; 14'h09F1: rddata <= 8'hAA; 14'h09F2: rddata <= 8'hBA; 14'h09F3: rddata <= 8'h57;
            14'h09F4: rddata <= 8'hDA; 14'h09F5: rddata <= 8'hC4; 14'h09F6: rddata <= 8'h03; 14'h09F7: rddata <= 8'h22;
            14'h09F8: rddata <= 8'hC3; 14'h09F9: rddata <= 8'h38; 14'h09FA: rddata <= 8'hD7; 14'h09FB: rddata <= 8'h18;
            14'h09FC: rddata <= 8'hE7; 14'h09FD: rddata <= 8'hF7; 14'h09FE: rddata <= 8'h09; 14'h09FF: rddata <= 8'hAF;
            14'h0A00: rddata <= 8'h32; 14'h0A01: rddata <= 8'hAB; 14'h0A02: rddata <= 8'h38; 14'h0A03: rddata <= 8'hD7;
            14'h0A04: rddata <= 8'hCA; 14'h0A05: rddata <= 8'hD6; 14'h0A06: rddata <= 8'h03; 14'h0A07: rddata <= 8'hDA;
            14'h0A08: rddata <= 8'hE5; 14'h0A09: rddata <= 8'h15; 14'h0A0A: rddata <= 8'hCD; 14'h0A0B: rddata <= 8'hC6;
            14'h0A0C: rddata <= 8'h0C; 14'h0A0D: rddata <= 8'hD2; 14'h0A0E: rddata <= 8'h4E; 14'h0A0F: rddata <= 8'h0A;
            14'h0A10: rddata <= 8'hFE; 14'h0A11: rddata <= 8'hA8; 14'h0A12: rddata <= 8'h28; 14'h0A13: rddata <= 8'hE9;
            14'h0A14: rddata <= 8'hFE; 14'h0A15: rddata <= 8'h2E; 14'h0A16: rddata <= 8'hCA; 14'h0A17: rddata <= 8'hE5;
            14'h0A18: rddata <= 8'h15; 14'h0A19: rddata <= 8'hFE; 14'h0A1A: rddata <= 8'hA9; 14'h0A1B: rddata <= 8'hCA;
            14'h0A1C: rddata <= 8'h3D; 14'h0A1D: rddata <= 8'h0A; 14'h0A1E: rddata <= 8'hFE; 14'h0A1F: rddata <= 8'h22;
            14'h0A20: rddata <= 8'hCA; 14'h0A21: rddata <= 8'h60; 14'h0A22: rddata <= 8'h0E; 14'h0A23: rddata <= 8'hFE;
            14'h0A24: rddata <= 8'hA6; 14'h0A25: rddata <= 8'hCA; 14'h0A26: rddata <= 8'h05; 14'h0A27: rddata <= 8'h0B;
            14'h0A28: rddata <= 8'hFE; 14'h0A29: rddata <= 8'hA4; 14'h0A2A: rddata <= 8'hCA; 14'h0A2B: rddata <= 8'hFB;
            14'h0A2C: rddata <= 8'h19; 14'h0A2D: rddata <= 8'hFE; 14'h0A2E: rddata <= 8'hA2; 14'h0A2F: rddata <= 8'hCA;
            14'h0A30: rddata <= 8'h40; 14'h0A31: rddata <= 8'h0B; 14'h0A32: rddata <= 8'hD6; 14'h0A33: rddata <= 8'hB2;
            14'h0A34: rddata <= 8'hD2; 14'h0A35: rddata <= 8'h5F; 14'h0A36: rddata <= 8'h0A; 14'h0A37: rddata <= 8'hCD;
            14'h0A38: rddata <= 8'h83; 14'h0A39: rddata <= 8'h09; 14'h0A3A: rddata <= 8'hCF; 14'h0A3B: rddata <= 8'h29;
            14'h0A3C: rddata <= 8'hC9; 14'h0A3D: rddata <= 8'h16; 14'h0A3E: rddata <= 8'h7D; 14'h0A3F: rddata <= 8'hCD;
            14'h0A40: rddata <= 8'h88; 14'h0A41: rddata <= 8'h09; 14'h0A42: rddata <= 8'h2A; 14'h0A43: rddata <= 8'hD0;
            14'h0A44: rddata <= 8'h38; 14'h0A45: rddata <= 8'hE5; 14'h0A46: rddata <= 8'hCD; 14'h0A47: rddata <= 8'h0B;
            14'h0A48: rddata <= 8'h15; 14'h0A49: rddata <= 8'hCD; 14'h0A4A: rddata <= 8'h75; 14'h0A4B: rddata <= 8'h09;
            14'h0A4C: rddata <= 8'hE1; 14'h0A4D: rddata <= 8'hC9; 14'h0A4E: rddata <= 8'hCD; 14'h0A4F: rddata <= 8'hD1;
            14'h0A50: rddata <= 8'h10; 14'h0A51: rddata <= 8'hE5; 14'h0A52: rddata <= 8'hEB; 14'h0A53: rddata <= 8'h22;
            14'h0A54: rddata <= 8'hE4; 14'h0A55: rddata <= 8'h38; 14'h0A56: rddata <= 8'h3A; 14'h0A57: rddata <= 8'hAB;
            14'h0A58: rddata <= 8'h38; 14'h0A59: rddata <= 8'hB7; 14'h0A5A: rddata <= 8'hCC; 14'h0A5B: rddata <= 8'h20;
            14'h0A5C: rddata <= 8'h15; 14'h0A5D: rddata <= 8'hE1; 14'h0A5E: rddata <= 8'hC9; 14'h0A5F: rddata <= 8'hF7;
            14'h0A60: rddata <= 8'h1B; 14'h0A61: rddata <= 8'hFE; 14'h0A62: rddata <= 8'h18; 14'h0A63: rddata <= 8'hCA;
            14'h0A64: rddata <= 8'h68; 14'h0A65: rddata <= 8'h1A; 14'h0A66: rddata <= 8'h06; 14'h0A67: rddata <= 8'h00;
            14'h0A68: rddata <= 8'h07; 14'h0A69: rddata <= 8'h4F; 14'h0A6A: rddata <= 8'hC5; 14'h0A6B: rddata <= 8'hD7;
            14'h0A6C: rddata <= 8'h79; 14'h0A6D: rddata <= 8'hFE; 14'h0A6E: rddata <= 8'h29; 14'h0A6F: rddata <= 8'h38;
            14'h0A70: rddata <= 8'h16; 14'h0A71: rddata <= 8'hCD; 14'h0A72: rddata <= 8'h83; 14'h0A73: rddata <= 8'h09;
            14'h0A74: rddata <= 8'hCF; 14'h0A75: rddata <= 8'h2C; 14'h0A76: rddata <= 8'hCD; 14'h0A77: rddata <= 8'h76;
            14'h0A78: rddata <= 8'h09; 14'h0A79: rddata <= 8'hEB; 14'h0A7A: rddata <= 8'h2A; 14'h0A7B: rddata <= 8'hE4;
            14'h0A7C: rddata <= 8'h38; 14'h0A7D: rddata <= 8'hE3; 14'h0A7E: rddata <= 8'hE5; 14'h0A7F: rddata <= 8'hEB;
            14'h0A80: rddata <= 8'hCD; 14'h0A81: rddata <= 8'h54; 14'h0A82: rddata <= 8'h0B; 14'h0A83: rddata <= 8'hEB;
            14'h0A84: rddata <= 8'hE3; 14'h0A85: rddata <= 8'h18; 14'h0A86: rddata <= 8'h08; 14'h0A87: rddata <= 8'hCD;
            14'h0A88: rddata <= 8'h37; 14'h0A89: rddata <= 8'h0A; 14'h0A8A: rddata <= 8'hE3; 14'h0A8B: rddata <= 8'h11;
            14'h0A8C: rddata <= 8'h49; 14'h0A8D: rddata <= 8'h0A; 14'h0A8E: rddata <= 8'hD5; 14'h0A8F: rddata <= 8'h01;
            14'h0A90: rddata <= 8'h15; 14'h0A91: rddata <= 8'h02; 14'h0A92: rddata <= 8'h09; 14'h0A93: rddata <= 8'h4E;
            14'h0A94: rddata <= 8'h23; 14'h0A95: rddata <= 8'h66; 14'h0A96: rddata <= 8'h69; 14'h0A97: rddata <= 8'hE9;
            14'h0A98: rddata <= 8'h15; 14'h0A99: rddata <= 8'hFE; 14'h0A9A: rddata <= 8'hA9; 14'h0A9B: rddata <= 8'hC8;
            14'h0A9C: rddata <= 8'hFE; 14'h0A9D: rddata <= 8'h2D; 14'h0A9E: rddata <= 8'hC8; 14'h0A9F: rddata <= 8'h14;
            14'h0AA0: rddata <= 8'hFE; 14'h0AA1: rddata <= 8'h2B; 14'h0AA2: rddata <= 8'hC8; 14'h0AA3: rddata <= 8'hFE;
            14'h0AA4: rddata <= 8'hA8; 14'h0AA5: rddata <= 8'hC8; 14'h0AA6: rddata <= 8'h2B; 14'h0AA7: rddata <= 8'hC9;
            14'h0AA8: rddata <= 8'hF6; 14'h0AA9: rddata <= 8'hAF; 14'h0AAA: rddata <= 8'hF5; 14'h0AAB: rddata <= 8'hCD;
            14'h0AAC: rddata <= 8'h75; 14'h0AAD: rddata <= 8'h09; 14'h0AAE: rddata <= 8'hCD; 14'h0AAF: rddata <= 8'h82;
            14'h0AB0: rddata <= 8'h06; 14'h0AB1: rddata <= 8'hF1; 14'h0AB2: rddata <= 8'hEB; 14'h0AB3: rddata <= 8'hC1;
            14'h0AB4: rddata <= 8'hE3; 14'h0AB5: rddata <= 8'hEB; 14'h0AB6: rddata <= 8'hCD; 14'h0AB7: rddata <= 8'h23;
            14'h0AB8: rddata <= 8'h15; 14'h0AB9: rddata <= 8'hF5; 14'h0ABA: rddata <= 8'hCD; 14'h0ABB: rddata <= 8'h82;
            14'h0ABC: rddata <= 8'h06; 14'h0ABD: rddata <= 8'hF1; 14'h0ABE: rddata <= 8'hC1; 14'h0ABF: rddata <= 8'h79;
            14'h0AC0: rddata <= 8'h21; 14'h0AC1: rddata <= 8'h21; 14'h0AC2: rddata <= 8'h0B; 14'h0AC3: rddata <= 8'hC2;
            14'h0AC4: rddata <= 8'hCB; 14'h0AC5: rddata <= 8'h0A; 14'h0AC6: rddata <= 8'hA3; 14'h0AC7: rddata <= 8'h4F;
            14'h0AC8: rddata <= 8'h78; 14'h0AC9: rddata <= 8'hA2; 14'h0ACA: rddata <= 8'hE9; 14'h0ACB: rddata <= 8'hB3;
            14'h0ACC: rddata <= 8'h4F; 14'h0ACD: rddata <= 8'h78; 14'h0ACE: rddata <= 8'hB2; 14'h0ACF: rddata <= 8'hE9;
            14'h0AD0: rddata <= 8'h21; 14'h0AD1: rddata <= 8'hE2; 14'h0AD2: rddata <= 8'h0A; 14'h0AD3: rddata <= 8'h3A;
            14'h0AD4: rddata <= 8'hAB; 14'h0AD5: rddata <= 8'h38; 14'h0AD6: rddata <= 8'h1F; 14'h0AD7: rddata <= 8'h7A;
            14'h0AD8: rddata <= 8'h17; 14'h0AD9: rddata <= 8'h5F; 14'h0ADA: rddata <= 8'h16; 14'h0ADB: rddata <= 8'h64;
            14'h0ADC: rddata <= 8'h78; 14'h0ADD: rddata <= 8'hBA; 14'h0ADE: rddata <= 8'hD0; 14'h0ADF: rddata <= 8'hC3;
            14'h0AE0: rddata <= 8'hCB; 14'h0AE1: rddata <= 8'h09; 14'h0AE2: rddata <= 8'hE4; 14'h0AE3: rddata <= 8'h0A;
            14'h0AE4: rddata <= 8'h79; 14'h0AE5: rddata <= 8'hB7; 14'h0AE6: rddata <= 8'h1F; 14'h0AE7: rddata <= 8'hC1;
            14'h0AE8: rddata <= 8'hD1; 14'h0AE9: rddata <= 8'hF5; 14'h0AEA: rddata <= 8'hCD; 14'h0AEB: rddata <= 8'h77;
            14'h0AEC: rddata <= 8'h09; 14'h0AED: rddata <= 8'h21; 14'h0AEE: rddata <= 8'hFB; 14'h0AEF: rddata <= 8'h0A;
            14'h0AF0: rddata <= 8'hE5; 14'h0AF1: rddata <= 8'hCA; 14'h0AF2: rddata <= 8'h5B; 14'h0AF3: rddata <= 8'h15;
            14'h0AF4: rddata <= 8'hAF; 14'h0AF5: rddata <= 8'h32; 14'h0AF6: rddata <= 8'hAB; 14'h0AF7: rddata <= 8'h38;
            14'h0AF8: rddata <= 8'hC3; 14'h0AF9: rddata <= 8'hFC; 14'h0AFA: rddata <= 8'h0D; 14'h0AFB: rddata <= 8'h3C;
            14'h0AFC: rddata <= 8'h8F; 14'h0AFD: rddata <= 8'hC1; 14'h0AFE: rddata <= 8'hA0; 14'h0AFF: rddata <= 8'hC6;
            14'h0B00: rddata <= 8'hFF; 14'h0B01: rddata <= 8'h9F; 14'h0B02: rddata <= 8'hC3; 14'h0B03: rddata <= 8'hF6;
            14'h0B04: rddata <= 8'h14; 14'h0B05: rddata <= 8'h16; 14'h0B06: rddata <= 8'h5A; 14'h0B07: rddata <= 8'hCD;
            14'h0B08: rddata <= 8'h88; 14'h0B09: rddata <= 8'h09; 14'h0B0A: rddata <= 8'hCD; 14'h0B0B: rddata <= 8'h75;
            14'h0B0C: rddata <= 8'h09; 14'h0B0D: rddata <= 8'hCD; 14'h0B0E: rddata <= 8'h82; 14'h0B0F: rddata <= 8'h06;
            14'h0B10: rddata <= 8'h7B; 14'h0B11: rddata <= 8'h2F; 14'h0B12: rddata <= 8'h4F; 14'h0B13: rddata <= 8'h7A;
            14'h0B14: rddata <= 8'h2F; 14'h0B15: rddata <= 8'hCD; 14'h0B16: rddata <= 8'h21; 14'h0B17: rddata <= 8'h0B;
            14'h0B18: rddata <= 8'hC1; 14'h0B19: rddata <= 8'hC3; 14'h0B1A: rddata <= 8'h94; 14'h0B1B: rddata <= 8'h09;
            14'h0B1C: rddata <= 8'h7D; 14'h0B1D: rddata <= 8'h93; 14'h0B1E: rddata <= 8'h4F; 14'h0B1F: rddata <= 8'h7C;
            14'h0B20: rddata <= 8'h9A; 14'h0B21: rddata <= 8'h41; 14'h0B22: rddata <= 8'h50; 14'h0B23: rddata <= 8'h1E;
            14'h0B24: rddata <= 8'h00; 14'h0B25: rddata <= 8'h21; 14'h0B26: rddata <= 8'hAB; 14'h0B27: rddata <= 8'h38;
            14'h0B28: rddata <= 8'h73; 14'h0B29: rddata <= 8'h06; 14'h0B2A: rddata <= 8'h90; 14'h0B2B: rddata <= 8'hC3;
            14'h0B2C: rddata <= 8'hFB; 14'h0B2D: rddata <= 8'h14; 14'h0B2E: rddata <= 8'h3A; 14'h0B2F: rddata <= 8'h46;
            14'h0B30: rddata <= 8'h38; 14'h0B31: rddata <= 8'h18; 14'h0B32: rddata <= 8'h03; 14'h0B33: rddata <= 8'h3A;
            14'h0B34: rddata <= 8'h00; 14'h0B35: rddata <= 8'h38; 14'h0B36: rddata <= 8'h47; 14'h0B37: rddata <= 8'hAF;
            14'h0B38: rddata <= 8'hC3; 14'h0B39: rddata <= 8'h22; 14'h0B3A: rddata <= 8'h0B; 14'h0B3B: rddata <= 8'hF7;
            14'h0B3C: rddata <= 8'h0F; 14'h0B3D: rddata <= 8'hC3; 14'h0B3E: rddata <= 8'hC4; 14'h0B3F: rddata <= 8'h03;
            14'h0B40: rddata <= 8'hF7; 14'h0B41: rddata <= 8'h10; 14'h0B42: rddata <= 8'hC3; 14'h0B43: rddata <= 8'hC4;
            14'h0B44: rddata <= 8'h03; 14'h0B45: rddata <= 8'hE5; 14'h0B46: rddata <= 8'h2A; 14'h0B47: rddata <= 8'h4D;
            14'h0B48: rddata <= 8'h38; 14'h0B49: rddata <= 8'h23; 14'h0B4A: rddata <= 8'h7C; 14'h0B4B: rddata <= 8'hB5;
            14'h0B4C: rddata <= 8'hE1; 14'h0B4D: rddata <= 8'hC0; 14'h0B4E: rddata <= 8'h1E; 14'h0B4F: rddata <= 8'h16;
            14'h0B50: rddata <= 8'hC3; 14'h0B51: rddata <= 8'hDB; 14'h0B52: rddata <= 8'h03; 14'h0B53: rddata <= 8'hD7;
            14'h0B54: rddata <= 8'hCD; 14'h0B55: rddata <= 8'h72; 14'h0B56: rddata <= 8'h09; 14'h0B57: rddata <= 8'hCD;
            14'h0B58: rddata <= 8'h7E; 14'h0B59: rddata <= 8'h06; 14'h0B5A: rddata <= 8'h7A; 14'h0B5B: rddata <= 8'hB7;
            14'h0B5C: rddata <= 8'hC2; 14'h0B5D: rddata <= 8'h97; 14'h0B5E: rddata <= 8'h06; 14'h0B5F: rddata <= 8'h2B;
            14'h0B60: rddata <= 8'hD7; 14'h0B61: rddata <= 8'h7B; 14'h0B62: rddata <= 8'hC9; 14'h0B63: rddata <= 8'hCD;
            14'h0B64: rddata <= 8'h82; 14'h0B65: rddata <= 8'h06; 14'h0B66: rddata <= 8'hCD; 14'h0B67: rddata <= 8'h88;
            14'h0B68: rddata <= 8'h0B; 14'h0B69: rddata <= 8'h1A; 14'h0B6A: rddata <= 8'hC3; 14'h0B6B: rddata <= 8'h36;
            14'h0B6C: rddata <= 8'h0B; 14'h0B6D: rddata <= 8'hCD; 14'h0B6E: rddata <= 8'h72; 14'h0B6F: rddata <= 8'h09;
            14'h0B70: rddata <= 8'hCD; 14'h0B71: rddata <= 8'h82; 14'h0B72: rddata <= 8'h06; 14'h0B73: rddata <= 8'hCD;
            14'h0B74: rddata <= 8'h88; 14'h0B75: rddata <= 8'h0B; 14'h0B76: rddata <= 8'hD5; 14'h0B77: rddata <= 8'hCF;
            14'h0B78: rddata <= 8'h2C; 14'h0B79: rddata <= 8'hCD; 14'h0B7A: rddata <= 8'h54; 14'h0B7B: rddata <= 8'h0B;
            14'h0B7C: rddata <= 8'hD1; 14'h0B7D: rddata <= 8'h12; 14'h0B7E: rddata <= 8'hC9; 14'h0B7F: rddata <= 8'hCD;
            14'h0B80: rddata <= 8'h85; 14'h0B81: rddata <= 8'h09; 14'h0B82: rddata <= 8'hE5; 14'h0B83: rddata <= 8'hCD;
            14'h0B84: rddata <= 8'h82; 14'h0B85: rddata <= 8'h06; 14'h0B86: rddata <= 8'hE1; 14'h0B87: rddata <= 8'hC9;
            14'h0B88: rddata <= 8'hE5; 14'h0B89: rddata <= 8'h21; 14'h0B8A: rddata <= 8'hFF; 14'h0B8B: rddata <= 8'h2F;
            14'h0B8C: rddata <= 8'hE7; 14'h0B8D: rddata <= 8'hE1; 14'h0B8E: rddata <= 8'hD2; 14'h0B8F: rddata <= 8'h97;
            14'h0B90: rddata <= 8'h06; 14'h0B91: rddata <= 8'hC9; 14'h0B92: rddata <= 8'hCD; 14'h0B93: rddata <= 8'hA9;
            14'h0B94: rddata <= 8'h0B; 14'h0B95: rddata <= 8'hC5; 14'h0B96: rddata <= 8'hE3; 14'h0B97: rddata <= 8'hC1;
            14'h0B98: rddata <= 8'hE7; 14'h0B99: rddata <= 8'h7E; 14'h0B9A: rddata <= 8'h02; 14'h0B9B: rddata <= 8'hC8;
            14'h0B9C: rddata <= 8'h0B; 14'h0B9D: rddata <= 8'h2B; 14'h0B9E: rddata <= 8'h18; 14'h0B9F: rddata <= 8'hF8;
            14'h0BA0: rddata <= 8'hE5; 14'h0BA1: rddata <= 8'h2A; 14'h0BA2: rddata <= 8'hDA; 14'h0BA3: rddata <= 8'h38;
            14'h0BA4: rddata <= 8'h06; 14'h0BA5: rddata <= 8'h00; 14'h0BA6: rddata <= 8'h09; 14'h0BA7: rddata <= 8'h09;
            14'h0BA8: rddata <= 8'h3E; 14'h0BA9: rddata <= 8'hE5; 14'h0BAA: rddata <= 8'h3E; 14'h0BAB: rddata <= 8'hD0;
            14'h0BAC: rddata <= 8'h95; 14'h0BAD: rddata <= 8'h6F; 14'h0BAE: rddata <= 8'h3E; 14'h0BAF: rddata <= 8'hFF;
            14'h0BB0: rddata <= 8'h9C; 14'h0BB1: rddata <= 8'h67; 14'h0BB2: rddata <= 8'h38; 14'h0BB3: rddata <= 8'h03;
            14'h0BB4: rddata <= 8'h39; 14'h0BB5: rddata <= 8'hE1; 14'h0BB6: rddata <= 8'hD8; 14'h0BB7: rddata <= 8'h11;
            14'h0BB8: rddata <= 8'h0C; 14'h0BB9: rddata <= 8'h00; 14'h0BBA: rddata <= 8'hC3; 14'h0BBB: rddata <= 8'hDB;
            14'h0BBC: rddata <= 8'h03; 14'h0BBD: rddata <= 8'hC0; 14'h0BBE: rddata <= 8'hF7; 14'h0BBF: rddata <= 8'h0C;
            14'h0BC0: rddata <= 8'h2A; 14'h0BC1: rddata <= 8'h4F; 14'h0BC2: rddata <= 8'h38; 14'h0BC3: rddata <= 8'hAF;
            14'h0BC4: rddata <= 8'h77; 14'h0BC5: rddata <= 8'h23; 14'h0BC6: rddata <= 8'h77; 14'h0BC7: rddata <= 8'h23;
            14'h0BC8: rddata <= 8'h22; 14'h0BC9: rddata <= 8'hD6; 14'h0BCA: rddata <= 8'h38; 14'h0BCB: rddata <= 8'h2A;
            14'h0BCC: rddata <= 8'h4F; 14'h0BCD: rddata <= 8'h38; 14'h0BCE: rddata <= 8'h2B; 14'h0BCF: rddata <= 8'h22;
            14'h0BD0: rddata <= 8'hCE; 14'h0BD1: rddata <= 8'h38; 14'h0BD2: rddata <= 8'h2A; 14'h0BD3: rddata <= 8'hAD;
            14'h0BD4: rddata <= 8'h38; 14'h0BD5: rddata <= 8'h22; 14'h0BD6: rddata <= 8'hC1; 14'h0BD7: rddata <= 8'h38;
            14'h0BD8: rddata <= 8'hAF; 14'h0BD9: rddata <= 8'hCD; 14'h0BDA: rddata <= 8'h05; 14'h0BDB: rddata <= 8'h0C;
            14'h0BDC: rddata <= 8'h2A; 14'h0BDD: rddata <= 8'hD6; 14'h0BDE: rddata <= 8'h38; 14'h0BDF: rddata <= 8'h22;
            14'h0BE0: rddata <= 8'hD8; 14'h0BE1: rddata <= 8'h38; 14'h0BE2: rddata <= 8'h22; 14'h0BE3: rddata <= 8'hDA;
            14'h0BE4: rddata <= 8'h38; 14'h0BE5: rddata <= 8'hC1; 14'h0BE6: rddata <= 8'h2A; 14'h0BE7: rddata <= 8'h4B;
            14'h0BE8: rddata <= 8'h38; 14'h0BE9: rddata <= 8'hF9; 14'h0BEA: rddata <= 8'hCD; 14'h0BEB: rddata <= 8'hD8;
            14'h0BEC: rddata <= 8'h1F; 14'h0BED: rddata <= 8'h22; 14'h0BEE: rddata <= 8'hAF; 14'h0BEF: rddata <= 8'h38;
            14'h0BF0: rddata <= 8'hCD; 14'h0BF1: rddata <= 8'hBE; 14'h0BF2: rddata <= 8'h19; 14'h0BF3: rddata <= 8'hAF;
            14'h0BF4: rddata <= 8'h6F; 14'h0BF5: rddata <= 8'h67; 14'h0BF6: rddata <= 8'h22; 14'h0BF7: rddata <= 8'hD4;
            14'h0BF8: rddata <= 8'h38; 14'h0BF9: rddata <= 8'h32; 14'h0BFA: rddata <= 8'hCB; 14'h0BFB: rddata <= 8'h38;
            14'h0BFC: rddata <= 8'h22; 14'h0BFD: rddata <= 8'hDE; 14'h0BFE: rddata <= 8'h38; 14'h0BFF: rddata <= 8'hE5;
            14'h0C00: rddata <= 8'hC5; 14'h0C01: rddata <= 8'h2A; 14'h0C02: rddata <= 8'hCE; 14'h0C03: rddata <= 8'h38;
            14'h0C04: rddata <= 8'hC9; 14'h0C05: rddata <= 8'hEB; 14'h0C06: rddata <= 8'h2A; 14'h0C07: rddata <= 8'h4F;
            14'h0C08: rddata <= 8'h38; 14'h0C09: rddata <= 8'h28; 14'h0C0A: rddata <= 8'h0E; 14'h0C0B: rddata <= 8'hEB;
            14'h0C0C: rddata <= 8'hCD; 14'h0C0D: rddata <= 8'h9C; 14'h0C0E: rddata <= 8'h06; 14'h0C0F: rddata <= 8'hE5;
            14'h0C10: rddata <= 8'hCD; 14'h0C11: rddata <= 8'h9F; 14'h0C12: rddata <= 8'h04; 14'h0C13: rddata <= 8'h60;
            14'h0C14: rddata <= 8'h69; 14'h0C15: rddata <= 8'hD1; 14'h0C16: rddata <= 8'hD2; 14'h0C17: rddata <= 8'hF3;
            14'h0C18: rddata <= 8'h06; 14'h0C19: rddata <= 8'h2B; 14'h0C1A: rddata <= 8'h22; 14'h0C1B: rddata <= 8'hDC;
            14'h0C1C: rddata <= 8'h38; 14'h0C1D: rddata <= 8'hEB; 14'h0C1E: rddata <= 8'hC9; 14'h0C1F: rddata <= 8'hC0;
            14'h0C20: rddata <= 8'hF6; 14'h0C21: rddata <= 8'hC0; 14'h0C22: rddata <= 8'h22; 14'h0C23: rddata <= 8'hCE;
            14'h0C24: rddata <= 8'h38; 14'h0C25: rddata <= 8'h21; 14'h0C26: rddata <= 8'hF6; 14'h0C27: rddata <= 8'hFF;
            14'h0C28: rddata <= 8'hC1; 14'h0C29: rddata <= 8'h2A; 14'h0C2A: rddata <= 8'h4D; 14'h0C2B: rddata <= 8'h38;
            14'h0C2C: rddata <= 8'hF5; 14'h0C2D: rddata <= 8'h7D; 14'h0C2E: rddata <= 8'hA4; 14'h0C2F: rddata <= 8'h3C;
            14'h0C30: rddata <= 8'h28; 14'h0C31: rddata <= 8'h09; 14'h0C32: rddata <= 8'h22; 14'h0C33: rddata <= 8'hD2;
            14'h0C34: rddata <= 8'h38; 14'h0C35: rddata <= 8'h2A; 14'h0C36: rddata <= 8'hCE; 14'h0C37: rddata <= 8'h38;
            14'h0C38: rddata <= 8'h22; 14'h0C39: rddata <= 8'hD4; 14'h0C3A: rddata <= 8'h38; 14'h0C3B: rddata <= 8'hCD;
            14'h0C3C: rddata <= 8'hBE; 14'h0C3D: rddata <= 8'h19; 14'h0C3E: rddata <= 8'hCD; 14'h0C3F: rddata <= 8'hDE;
            14'h0C40: rddata <= 8'h19; 14'h0C41: rddata <= 8'hF1; 14'h0C42: rddata <= 8'h21; 14'h0C43: rddata <= 8'h73;
            14'h0C44: rddata <= 8'h03; 14'h0C45: rddata <= 8'hC2; 14'h0C46: rddata <= 8'hF4; 14'h0C47: rddata <= 8'h03;
            14'h0C48: rddata <= 8'hC3; 14'h0C49: rddata <= 8'h02; 14'h0C4A: rddata <= 8'h04; 14'h0C4B: rddata <= 8'h2A;
            14'h0C4C: rddata <= 8'hD4; 14'h0C4D: rddata <= 8'h38; 14'h0C4E: rddata <= 8'h7C; 14'h0C4F: rddata <= 8'hB5;
            14'h0C50: rddata <= 8'h11; 14'h0C51: rddata <= 8'h20; 14'h0C52: rddata <= 8'h00; 14'h0C53: rddata <= 8'hCA;
            14'h0C54: rddata <= 8'hDB; 14'h0C55: rddata <= 8'h03; 14'h0C56: rddata <= 8'hED; 14'h0C57: rddata <= 8'h5B;
            14'h0C58: rddata <= 8'hD2; 14'h0C59: rddata <= 8'h38; 14'h0C5A: rddata <= 8'hED; 14'h0C5B: rddata <= 8'h53;
            14'h0C5C: rddata <= 8'h4D; 14'h0C5D: rddata <= 8'h38; 14'h0C5E: rddata <= 8'hC9; 14'h0C5F: rddata <= 8'hC3;
            14'h0C60: rddata <= 8'h97; 14'h0C61: rddata <= 8'h06; 14'h0C62: rddata <= 8'h3E; 14'h0C63: rddata <= 8'hAF;
            14'h0C64: rddata <= 8'hB7; 14'h0C65: rddata <= 8'hF5; 14'h0C66: rddata <= 8'hD7; 14'h0C67: rddata <= 8'h3E;
            14'h0C68: rddata <= 8'h01; 14'h0C69: rddata <= 8'h32; 14'h0C6A: rddata <= 8'hCB; 14'h0C6B: rddata <= 8'h38;
            14'h0C6C: rddata <= 8'hCD; 14'h0C6D: rddata <= 8'hD1; 14'h0C6E: rddata <= 8'h10; 14'h0C6F: rddata <= 8'hC2;
            14'h0C70: rddata <= 8'h97; 14'h0C71: rddata <= 8'h06; 14'h0C72: rddata <= 8'h32; 14'h0C73: rddata <= 8'hCB;
            14'h0C74: rddata <= 8'h38; 14'h0C75: rddata <= 8'hCD; 14'h0C76: rddata <= 8'h75; 14'h0C77: rddata <= 8'h09;
            14'h0C78: rddata <= 8'hF1; 14'h0C79: rddata <= 8'hE5; 14'h0C7A: rddata <= 8'hF5; 14'h0C7B: rddata <= 8'hC5;
            14'h0C7C: rddata <= 8'h06; 14'h0C7D: rddata <= 8'h23; 14'h0C7E: rddata <= 8'h28; 14'h0C7F: rddata <= 8'h12;
            14'h0C80: rddata <= 8'hCD; 14'h0C81: rddata <= 8'h7F; 14'h0C82: rddata <= 8'h1B; 14'h0C83: rddata <= 8'hCD;
            14'h0C84: rddata <= 8'hBC; 14'h0C85: rddata <= 8'h1B; 14'h0C86: rddata <= 8'h78; 14'h0C87: rddata <= 8'hCD;
            14'h0C88: rddata <= 8'h87; 14'h0C89: rddata <= 8'h1B; 14'h0C8A: rddata <= 8'hCD; 14'h0C8B: rddata <= 8'h87;
            14'h0C8C: rddata <= 8'h1B; 14'h0C8D: rddata <= 8'hCD; 14'h0C8E: rddata <= 8'h87; 14'h0C8F: rddata <= 8'h1B;
            14'h0C90: rddata <= 8'h18; 14'h0C91: rddata <= 8'h11; 14'h0C92: rddata <= 8'hCD; 14'h0C93: rddata <= 8'h2E;
            14'h0C94: rddata <= 8'h1B; 14'h0C95: rddata <= 8'hCD; 14'h0C96: rddata <= 8'hCE; 14'h0C97: rddata <= 8'h1B;
            14'h0C98: rddata <= 8'h0E; 14'h0C99: rddata <= 8'h06; 14'h0C9A: rddata <= 8'hCD; 14'h0C9B: rddata <= 8'h4D;
            14'h0C9C: rddata <= 8'h1B; 14'h0C9D: rddata <= 8'hB8; 14'h0C9E: rddata <= 8'h20; 14'h0C9F: rddata <= 8'hF8;
            14'h0CA0: rddata <= 8'h0D; 14'h0CA1: rddata <= 8'h20; 14'h0CA2: rddata <= 8'hF7; 14'h0CA3: rddata <= 8'hE1;
            14'h0CA4: rddata <= 8'hEB; 14'h0CA5: rddata <= 8'h19; 14'h0CA6: rddata <= 8'hEB; 14'h0CA7: rddata <= 8'h4E;
            14'h0CA8: rddata <= 8'h06; 14'h0CA9: rddata <= 8'h00; 14'h0CAA: rddata <= 8'h09; 14'h0CAB: rddata <= 8'h09;
            14'h0CAC: rddata <= 8'h23; 14'h0CAD: rddata <= 8'hE7; 14'h0CAE: rddata <= 8'h28; 14'h0CAF: rddata <= 8'h0D;
            14'h0CB0: rddata <= 8'hF1; 14'h0CB1: rddata <= 8'hF5; 14'h0CB2: rddata <= 8'h7E; 14'h0CB3: rddata <= 8'hC4;
            14'h0CB4: rddata <= 8'h8A; 14'h0CB5: rddata <= 8'h1B; 14'h0CB6: rddata <= 8'hCC; 14'h0CB7: rddata <= 8'h4D;
            14'h0CB8: rddata <= 8'h1B; 14'h0CB9: rddata <= 8'h77; 14'h0CBA: rddata <= 8'h23; 14'h0CBB: rddata <= 8'h18;
            14'h0CBC: rddata <= 8'hF0; 14'h0CBD: rddata <= 8'hF1; 14'h0CBE: rddata <= 8'hC2; 14'h0CBF: rddata <= 8'h1C;
            14'h0CC0: rddata <= 8'h1C; 14'h0CC1: rddata <= 8'hE1; 14'h0CC2: rddata <= 8'hC3; 14'h0CC3: rddata <= 8'h7E;
            14'h0CC4: rddata <= 8'h1B; 14'h0CC5: rddata <= 8'h7E; 14'h0CC6: rddata <= 8'hFE; 14'h0CC7: rddata <= 8'h41;
            14'h0CC8: rddata <= 8'hD8; 14'h0CC9: rddata <= 8'hFE; 14'h0CCA: rddata <= 8'h5B; 14'h0CCB: rddata <= 8'h3F;
            14'h0CCC: rddata <= 8'hC9; 14'h0CCD: rddata <= 8'hF7; 14'h0CCE: rddata <= 8'h0B; 14'h0CCF: rddata <= 8'hCA;
            14'h0CD0: rddata <= 8'hCF; 14'h0CD1: rddata <= 8'h0B; 14'h0CD2: rddata <= 8'hCD; 14'h0CD3: rddata <= 8'h7B;
            14'h0CD4: rddata <= 8'h06; 14'h0CD5: rddata <= 8'h2B; 14'h0CD6: rddata <= 8'hD7; 14'h0CD7: rddata <= 8'hE5;
            14'h0CD8: rddata <= 8'h2A; 14'h0CD9: rddata <= 8'hAD; 14'h0CDA: rddata <= 8'h38; 14'h0CDB: rddata <= 8'h28;
            14'h0CDC: rddata <= 8'h0E; 14'h0CDD: rddata <= 8'hE1; 14'h0CDE: rddata <= 8'hCF; 14'h0CDF: rddata <= 8'h2C;
            14'h0CE0: rddata <= 8'hD5; 14'h0CE1: rddata <= 8'hCD; 14'h0CE2: rddata <= 8'h7B; 14'h0CE3: rddata <= 8'h06;
            14'h0CE4: rddata <= 8'h2B; 14'h0CE5: rddata <= 8'hD7; 14'h0CE6: rddata <= 8'hC2; 14'h0CE7: rddata <= 8'hC4;
            14'h0CE8: rddata <= 8'h03; 14'h0CE9: rddata <= 8'hE3; 14'h0CEA: rddata <= 8'hEB; 14'h0CEB: rddata <= 8'h7D;
            14'h0CEC: rddata <= 8'h93; 14'h0CED: rddata <= 8'h5F; 14'h0CEE: rddata <= 8'h7C; 14'h0CEF: rddata <= 8'h9A;
            14'h0CF0: rddata <= 8'h57; 14'h0CF1: rddata <= 8'hDA; 14'h0CF2: rddata <= 8'hB7; 14'h0CF3: rddata <= 8'h0B;
            14'h0CF4: rddata <= 8'hE5; 14'h0CF5: rddata <= 8'h2A; 14'h0CF6: rddata <= 8'hD6; 14'h0CF7: rddata <= 8'h38;
            14'h0CF8: rddata <= 8'h01; 14'h0CF9: rddata <= 8'h28; 14'h0CFA: rddata <= 8'h00; 14'h0CFB: rddata <= 8'h09;
            14'h0CFC: rddata <= 8'hE7; 14'h0CFD: rddata <= 8'hD2; 14'h0CFE: rddata <= 8'hB7; 14'h0CFF: rddata <= 8'h0B;
            14'h0D00: rddata <= 8'hEB; 14'h0D01: rddata <= 8'h22; 14'h0D02: rddata <= 8'h4B; 14'h0D03: rddata <= 8'h38;
            14'h0D04: rddata <= 8'hE1; 14'h0D05: rddata <= 8'h22; 14'h0D06: rddata <= 8'hAD; 14'h0D07: rddata <= 8'h38;
            14'h0D08: rddata <= 8'hE1; 14'h0D09: rddata <= 8'hC3; 14'h0D0A: rddata <= 8'hCF; 14'h0D0B: rddata <= 8'h0B;
            14'h0D0C: rddata <= 8'h7D; 14'h0D0D: rddata <= 8'h93; 14'h0D0E: rddata <= 8'h5F; 14'h0D0F: rddata <= 8'h7C;
            14'h0D10: rddata <= 8'h9A; 14'h0D11: rddata <= 8'h57; 14'h0D12: rddata <= 8'hC9; 14'h0D13: rddata <= 8'h11;
            14'h0D14: rddata <= 8'h00; 14'h0D15: rddata <= 8'h00; 14'h0D16: rddata <= 8'hC4; 14'h0D17: rddata <= 8'hD1;
            14'h0D18: rddata <= 8'h10; 14'h0D19: rddata <= 8'h22; 14'h0D1A: rddata <= 8'hCE; 14'h0D1B: rddata <= 8'h38;
            14'h0D1C: rddata <= 8'hCD; 14'h0D1D: rddata <= 8'h9F; 14'h0D1E: rddata <= 8'h03; 14'h0D1F: rddata <= 8'hC2;
            14'h0D20: rddata <= 8'hCA; 14'h0D21: rddata <= 8'h03; 14'h0D22: rddata <= 8'hF9; 14'h0D23: rddata <= 8'hD5;
            14'h0D24: rddata <= 8'h7E; 14'h0D25: rddata <= 8'hF5; 14'h0D26: rddata <= 8'h23; 14'h0D27: rddata <= 8'hD5;
            14'h0D28: rddata <= 8'hCD; 14'h0D29: rddata <= 8'h20; 14'h0D2A: rddata <= 8'h15; 14'h0D2B: rddata <= 8'hE3;
            14'h0D2C: rddata <= 8'hE5; 14'h0D2D: rddata <= 8'hCD; 14'h0D2E: rddata <= 8'h53; 14'h0D2F: rddata <= 8'h12;
            14'h0D30: rddata <= 8'hE1; 14'h0D31: rddata <= 8'hCD; 14'h0D32: rddata <= 8'h3A; 14'h0D33: rddata <= 8'h15;
            14'h0D34: rddata <= 8'hE1; 14'h0D35: rddata <= 8'hCD; 14'h0D36: rddata <= 8'h31; 14'h0D37: rddata <= 8'h15;
            14'h0D38: rddata <= 8'hE5; 14'h0D39: rddata <= 8'hCD; 14'h0D3A: rddata <= 8'h5B; 14'h0D3B: rddata <= 8'h15;
            14'h0D3C: rddata <= 8'hE1; 14'h0D3D: rddata <= 8'hC1; 14'h0D3E: rddata <= 8'h90; 14'h0D3F: rddata <= 8'hCD;
            14'h0D40: rddata <= 8'h31; 14'h0D41: rddata <= 8'h15; 14'h0D42: rddata <= 8'h28; 14'h0D43: rddata <= 8'h09;
            14'h0D44: rddata <= 8'hEB; 14'h0D45: rddata <= 8'h22; 14'h0D46: rddata <= 8'h4D; 14'h0D47: rddata <= 8'h38;
            14'h0D48: rddata <= 8'h69; 14'h0D49: rddata <= 8'h60; 14'h0D4A: rddata <= 8'hC3; 14'h0D4B: rddata <= 8'h28;
            14'h0D4C: rddata <= 8'h06; 14'h0D4D: rddata <= 8'hF9; 14'h0D4E: rddata <= 8'h2A; 14'h0D4F: rddata <= 8'hCE;
            14'h0D50: rddata <= 8'h38; 14'h0D51: rddata <= 8'h7E; 14'h0D52: rddata <= 8'hFE; 14'h0D53: rddata <= 8'h2C;
            14'h0D54: rddata <= 8'hC2; 14'h0D55: rddata <= 8'h2C; 14'h0D56: rddata <= 8'h06; 14'h0D57: rddata <= 8'hD7;
            14'h0D58: rddata <= 8'hCD; 14'h0D59: rddata <= 8'h16; 14'h0D5A: rddata <= 8'h0D; 14'h0D5B: rddata <= 8'h3E;
            14'h0D5C: rddata <= 8'h3F; 14'h0D5D: rddata <= 8'hDF; 14'h0D5E: rddata <= 8'h3E; 14'h0D5F: rddata <= 8'h20;
            14'h0D60: rddata <= 8'hDF; 14'h0D61: rddata <= 8'hC3; 14'h0D62: rddata <= 8'h85; 14'h0D63: rddata <= 8'h0D;
            14'h0D64: rddata <= 8'h3A; 14'h0D65: rddata <= 8'h4A; 14'h0D66: rddata <= 8'h38; 14'h0D67: rddata <= 8'hB7;
            14'h0D68: rddata <= 8'h3E; 14'h0D69: rddata <= 8'h5C; 14'h0D6A: rddata <= 8'h32; 14'h0D6B: rddata <= 8'h4A;
            14'h0D6C: rddata <= 8'h38; 14'h0D6D: rddata <= 8'h20; 14'h0D6E: rddata <= 8'h05; 14'h0D6F: rddata <= 8'h05;
            14'h0D70: rddata <= 8'h28; 14'h0D71: rddata <= 8'h13; 14'h0D72: rddata <= 8'hDF; 14'h0D73: rddata <= 8'h04;
            14'h0D74: rddata <= 8'h05; 14'h0D75: rddata <= 8'h2B; 14'h0D76: rddata <= 8'h28; 14'h0D77: rddata <= 8'h09;
            14'h0D78: rddata <= 8'h7E; 14'h0D79: rddata <= 8'hDF; 14'h0D7A: rddata <= 8'h18; 14'h0D7B: rddata <= 8'h12;
            14'h0D7C: rddata <= 8'h05; 14'h0D7D: rddata <= 8'h2B; 14'h0D7E: rddata <= 8'hDF; 14'h0D7F: rddata <= 8'h20;
            14'h0D80: rddata <= 8'h0D; 14'h0D81: rddata <= 8'hDF; 14'h0D82: rddata <= 8'hCD; 14'h0D83: rddata <= 8'hEA;
            14'h0D84: rddata <= 8'h19; 14'h0D85: rddata <= 8'h21; 14'h0D86: rddata <= 8'h60; 14'h0D87: rddata <= 8'h38;
            14'h0D88: rddata <= 8'h06; 14'h0D89: rddata <= 8'h01; 14'h0D8A: rddata <= 8'hAF; 14'h0D8B: rddata <= 8'h32;
            14'h0D8C: rddata <= 8'h4A; 14'h0D8D: rddata <= 8'h38; 14'h0D8E: rddata <= 8'hCD; 14'h0D8F: rddata <= 8'hDA;
            14'h0D90: rddata <= 8'h19; 14'h0D91: rddata <= 8'h4F; 14'h0D92: rddata <= 8'hFE; 14'h0D93: rddata <= 8'h7F;
            14'h0D94: rddata <= 8'h28; 14'h0D95: rddata <= 8'hCE; 14'h0D96: rddata <= 8'h3A; 14'h0D97: rddata <= 8'h4A;
            14'h0D98: rddata <= 8'h38; 14'h0D99: rddata <= 8'hB7; 14'h0D9A: rddata <= 8'h28; 14'h0D9B: rddata <= 8'h07;
            14'h0D9C: rddata <= 8'h3E; 14'h0D9D: rddata <= 8'h5C; 14'h0D9E: rddata <= 8'hDF; 14'h0D9F: rddata <= 8'hAF;
            14'h0DA0: rddata <= 8'h32; 14'h0DA1: rddata <= 8'h4A; 14'h0DA2: rddata <= 8'h38; 14'h0DA3: rddata <= 8'h79;
            14'h0DA4: rddata <= 8'hFE; 14'h0DA5: rddata <= 8'h07; 14'h0DA6: rddata <= 8'h28; 14'h0DA7: rddata <= 8'h41;
            14'h0DA8: rddata <= 8'hFE; 14'h0DA9: rddata <= 8'h03; 14'h0DAA: rddata <= 8'hCC; 14'h0DAB: rddata <= 8'hEA;
            14'h0DAC: rddata <= 8'h19; 14'h0DAD: rddata <= 8'h37; 14'h0DAE: rddata <= 8'hC8; 14'h0DAF: rddata <= 8'hFE;
            14'h0DB0: rddata <= 8'h0D; 14'h0DB1: rddata <= 8'hCA; 14'h0DB2: rddata <= 8'hE5; 14'h0DB3: rddata <= 8'h19;
            14'h0DB4: rddata <= 8'hFE; 14'h0DB5: rddata <= 8'h15; 14'h0DB6: rddata <= 8'hCA; 14'h0DB7: rddata <= 8'h82;
            14'h0DB8: rddata <= 8'h0D; 14'h0DB9: rddata <= 8'h00; 14'h0DBA: rddata <= 8'h00; 14'h0DBB: rddata <= 8'h00;
            14'h0DBC: rddata <= 8'h00; 14'h0DBD: rddata <= 8'h00; 14'h0DBE: rddata <= 8'hFE; 14'h0DBF: rddata <= 8'h08;
            14'h0DC0: rddata <= 8'hCA; 14'h0DC1: rddata <= 8'h7C; 14'h0DC2: rddata <= 8'h0D; 14'h0DC3: rddata <= 8'hFE;
            14'h0DC4: rddata <= 8'h18; 14'h0DC5: rddata <= 8'h20; 14'h0DC6: rddata <= 8'h05; 14'h0DC7: rddata <= 8'h3E;
            14'h0DC8: rddata <= 8'h23; 14'h0DC9: rddata <= 8'hC3; 14'h0DCA: rddata <= 8'h81; 14'h0DCB: rddata <= 8'h0D;
            14'h0DCC: rddata <= 8'hFE; 14'h0DCD: rddata <= 8'h12; 14'h0DCE: rddata <= 8'h20; 14'h0DCF: rddata <= 8'h14;
            14'h0DD0: rddata <= 8'hC5; 14'h0DD1: rddata <= 8'hD5; 14'h0DD2: rddata <= 8'hE5; 14'h0DD3: rddata <= 8'h36;
            14'h0DD4: rddata <= 8'h00; 14'h0DD5: rddata <= 8'hCD; 14'h0DD6: rddata <= 8'hEA; 14'h0DD7: rddata <= 8'h19;
            14'h0DD8: rddata <= 8'h21; 14'h0DD9: rddata <= 8'h60; 14'h0DDA: rddata <= 8'h38; 14'h0DDB: rddata <= 8'hCD;
            14'h0DDC: rddata <= 8'h9D; 14'h0DDD: rddata <= 8'h0E; 14'h0DDE: rddata <= 8'hE1; 14'h0DDF: rddata <= 8'hD1;
            14'h0DE0: rddata <= 8'hC1; 14'h0DE1: rddata <= 8'hC3; 14'h0DE2: rddata <= 8'h8E; 14'h0DE3: rddata <= 8'h0D;
            14'h0DE4: rddata <= 8'hFE; 14'h0DE5: rddata <= 8'h20; 14'h0DE6: rddata <= 8'hDA; 14'h0DE7: rddata <= 8'h8E;
            14'h0DE8: rddata <= 8'h0D; 14'h0DE9: rddata <= 8'h78; 14'h0DEA: rddata <= 8'hFE; 14'h0DEB: rddata <= 8'h49;
            14'h0DEC: rddata <= 8'h3E; 14'h0DED: rddata <= 8'h07; 14'h0DEE: rddata <= 8'hD2; 14'h0DEF: rddata <= 8'hF8;
            14'h0DF0: rddata <= 8'h0D; 14'h0DF1: rddata <= 8'h79; 14'h0DF2: rddata <= 8'h71; 14'h0DF3: rddata <= 8'h32;
            14'h0DF4: rddata <= 8'hCC; 14'h0DF5: rddata <= 8'h38; 14'h0DF6: rddata <= 8'h23; 14'h0DF7: rddata <= 8'h04;
            14'h0DF8: rddata <= 8'hDF; 14'h0DF9: rddata <= 8'hC3; 14'h0DFA: rddata <= 8'h8E; 14'h0DFB: rddata <= 8'h0D;
            14'h0DFC: rddata <= 8'hD5; 14'h0DFD: rddata <= 8'hCD; 14'h0DFE: rddata <= 8'hC9; 14'h0DFF: rddata <= 8'h0F;
            14'h0E00: rddata <= 8'h7E; 14'h0E01: rddata <= 8'h23; 14'h0E02: rddata <= 8'h23; 14'h0E03: rddata <= 8'h4E;
            14'h0E04: rddata <= 8'h23; 14'h0E05: rddata <= 8'h46; 14'h0E06: rddata <= 8'hD1; 14'h0E07: rddata <= 8'hC5;
            14'h0E08: rddata <= 8'hF5; 14'h0E09: rddata <= 8'hCD; 14'h0E0A: rddata <= 8'hCD; 14'h0E0B: rddata <= 8'h0F;
            14'h0E0C: rddata <= 8'hCD; 14'h0E0D: rddata <= 8'h31; 14'h0E0E: rddata <= 8'h15; 14'h0E0F: rddata <= 8'hF1;
            14'h0E10: rddata <= 8'h57; 14'h0E11: rddata <= 8'hE1; 14'h0E12: rddata <= 8'h7B; 14'h0E13: rddata <= 8'hB2;
            14'h0E14: rddata <= 8'hC8; 14'h0E15: rddata <= 8'h7A; 14'h0E16: rddata <= 8'hD6; 14'h0E17: rddata <= 8'h01;
            14'h0E18: rddata <= 8'hD8; 14'h0E19: rddata <= 8'hAF; 14'h0E1A: rddata <= 8'hBB; 14'h0E1B: rddata <= 8'h3C;
            14'h0E1C: rddata <= 8'hD0; 14'h0E1D: rddata <= 8'h15; 14'h0E1E: rddata <= 8'h1D; 14'h0E1F: rddata <= 8'h0A;
            14'h0E20: rddata <= 8'h03; 14'h0E21: rddata <= 8'hBE; 14'h0E22: rddata <= 8'h23; 14'h0E23: rddata <= 8'h28;
            14'h0E24: rddata <= 8'hED; 14'h0E25: rddata <= 8'h3F; 14'h0E26: rddata <= 8'hC3; 14'h0E27: rddata <= 8'hF1;
            14'h0E28: rddata <= 8'h14; 14'h0E29: rddata <= 8'hCD; 14'h0E2A: rddata <= 8'h75; 14'h0E2B: rddata <= 8'h09;
            14'h0E2C: rddata <= 8'hCD; 14'h0E2D: rddata <= 8'h80; 14'h0E2E: rddata <= 8'h16; 14'h0E2F: rddata <= 8'hCD;
            14'h0E30: rddata <= 8'h5F; 14'h0E31: rddata <= 8'h0E; 14'h0E32: rddata <= 8'hCD; 14'h0E33: rddata <= 8'hC9;
            14'h0E34: rddata <= 8'h0F; 14'h0E35: rddata <= 8'h01; 14'h0E36: rddata <= 8'h1D; 14'h0E37: rddata <= 8'h10;
            14'h0E38: rddata <= 8'hC5; 14'h0E39: rddata <= 8'h7E; 14'h0E3A: rddata <= 8'h23; 14'h0E3B: rddata <= 8'h23;
            14'h0E3C: rddata <= 8'hE5; 14'h0E3D: rddata <= 8'hCD; 14'h0E3E: rddata <= 8'hB3; 14'h0E3F: rddata <= 8'h0E;
            14'h0E40: rddata <= 8'hE1; 14'h0E41: rddata <= 8'h4E; 14'h0E42: rddata <= 8'h23; 14'h0E43: rddata <= 8'h46;
            14'h0E44: rddata <= 8'hCD; 14'h0E45: rddata <= 8'h53; 14'h0E46: rddata <= 8'h0E; 14'h0E47: rddata <= 8'hE5;
            14'h0E48: rddata <= 8'h6F; 14'h0E49: rddata <= 8'hCD; 14'h0E4A: rddata <= 8'hBD; 14'h0E4B: rddata <= 8'h0F;
            14'h0E4C: rddata <= 8'hD1; 14'h0E4D: rddata <= 8'hC9; 14'h0E4E: rddata <= 8'h3E; 14'h0E4F: rddata <= 8'h01;
            14'h0E50: rddata <= 8'hCD; 14'h0E51: rddata <= 8'hB3; 14'h0E52: rddata <= 8'h0E; 14'h0E53: rddata <= 8'h21;
            14'h0E54: rddata <= 8'hBD; 14'h0E55: rddata <= 8'h38; 14'h0E56: rddata <= 8'hE5; 14'h0E57: rddata <= 8'h77;
            14'h0E58: rddata <= 8'h23; 14'h0E59: rddata <= 8'h23; 14'h0E5A: rddata <= 8'h73; 14'h0E5B: rddata <= 8'h23;
            14'h0E5C: rddata <= 8'h72; 14'h0E5D: rddata <= 8'hE1; 14'h0E5E: rddata <= 8'hC9; 14'h0E5F: rddata <= 8'h2B;
            14'h0E60: rddata <= 8'h06; 14'h0E61: rddata <= 8'h22; 14'h0E62: rddata <= 8'h50; 14'h0E63: rddata <= 8'hE5;
            14'h0E64: rddata <= 8'h0E; 14'h0E65: rddata <= 8'hFF; 14'h0E66: rddata <= 8'h23; 14'h0E67: rddata <= 8'h7E;
            14'h0E68: rddata <= 8'h0C; 14'h0E69: rddata <= 8'hB7; 14'h0E6A: rddata <= 8'h28; 14'h0E6B: rddata <= 8'h06;
            14'h0E6C: rddata <= 8'hBA; 14'h0E6D: rddata <= 8'h28; 14'h0E6E: rddata <= 8'h03; 14'h0E6F: rddata <= 8'hB8;
            14'h0E70: rddata <= 8'h20; 14'h0E71: rddata <= 8'hF4; 14'h0E72: rddata <= 8'hFE; 14'h0E73: rddata <= 8'h22;
            14'h0E74: rddata <= 8'hCC; 14'h0E75: rddata <= 8'h6B; 14'h0E76: rddata <= 8'h06; 14'h0E77: rddata <= 8'hE3;
            14'h0E78: rddata <= 8'h23; 14'h0E79: rddata <= 8'hEB; 14'h0E7A: rddata <= 8'h79; 14'h0E7B: rddata <= 8'hCD;
            14'h0E7C: rddata <= 8'h53; 14'h0E7D: rddata <= 8'h0E; 14'h0E7E: rddata <= 8'h11; 14'h0E7F: rddata <= 8'hBD;
            14'h0E80: rddata <= 8'h38; 14'h0E81: rddata <= 8'h2A; 14'h0E82: rddata <= 8'hAF; 14'h0E83: rddata <= 8'h38;
            14'h0E84: rddata <= 8'h22; 14'h0E85: rddata <= 8'hE4; 14'h0E86: rddata <= 8'h38; 14'h0E87: rddata <= 8'h3E;
            14'h0E88: rddata <= 8'h01; 14'h0E89: rddata <= 8'h32; 14'h0E8A: rddata <= 8'hAB; 14'h0E8B: rddata <= 8'h38;
            14'h0E8C: rddata <= 8'hCD; 14'h0E8D: rddata <= 8'h3D; 14'h0E8E: rddata <= 8'h15; 14'h0E8F: rddata <= 8'hE7;
            14'h0E90: rddata <= 8'h22; 14'h0E91: rddata <= 8'hAF; 14'h0E92: rddata <= 8'h38; 14'h0E93: rddata <= 8'hE1;
            14'h0E94: rddata <= 8'h7E; 14'h0E95: rddata <= 8'hC0; 14'h0E96: rddata <= 8'h11; 14'h0E97: rddata <= 8'h1E;
            14'h0E98: rddata <= 8'h00; 14'h0E99: rddata <= 8'hC3; 14'h0E9A: rddata <= 8'hDB; 14'h0E9B: rddata <= 8'h03;
            14'h0E9C: rddata <= 8'h23; 14'h0E9D: rddata <= 8'hCD; 14'h0E9E: rddata <= 8'h5F; 14'h0E9F: rddata <= 8'h0E;
            14'h0EA0: rddata <= 8'hCD; 14'h0EA1: rddata <= 8'hC9; 14'h0EA2: rddata <= 8'h0F; 14'h0EA3: rddata <= 8'hCD;
            14'h0EA4: rddata <= 8'h31; 14'h0EA5: rddata <= 8'h15; 14'h0EA6: rddata <= 8'h1C; 14'h0EA7: rddata <= 8'h1D;
            14'h0EA8: rddata <= 8'hC8; 14'h0EA9: rddata <= 8'h0A; 14'h0EAA: rddata <= 8'hDF; 14'h0EAB: rddata <= 8'hFE;
            14'h0EAC: rddata <= 8'h0D; 14'h0EAD: rddata <= 8'hCC; 14'h0EAE: rddata <= 8'hF0; 14'h0EAF: rddata <= 8'h19;
            14'h0EB0: rddata <= 8'h03; 14'h0EB1: rddata <= 8'h18; 14'h0EB2: rddata <= 8'hF4; 14'h0EB3: rddata <= 8'hB7;
            14'h0EB4: rddata <= 8'h0E; 14'h0EB5: rddata <= 8'hF1; 14'h0EB6: rddata <= 8'hF5; 14'h0EB7: rddata <= 8'h2A;
            14'h0EB8: rddata <= 8'h4B; 14'h0EB9: rddata <= 8'h38; 14'h0EBA: rddata <= 8'hEB; 14'h0EBB: rddata <= 8'h2A;
            14'h0EBC: rddata <= 8'hC1; 14'h0EBD: rddata <= 8'h38; 14'h0EBE: rddata <= 8'h2F; 14'h0EBF: rddata <= 8'h4F;
            14'h0EC0: rddata <= 8'h06; 14'h0EC1: rddata <= 8'hFF; 14'h0EC2: rddata <= 8'h09; 14'h0EC3: rddata <= 8'h23;
            14'h0EC4: rddata <= 8'hE7; 14'h0EC5: rddata <= 8'h38; 14'h0EC6: rddata <= 8'h07; 14'h0EC7: rddata <= 8'h22;
            14'h0EC8: rddata <= 8'hC1; 14'h0EC9: rddata <= 8'h38; 14'h0ECA: rddata <= 8'h23; 14'h0ECB: rddata <= 8'hEB;
            14'h0ECC: rddata <= 8'hF1; 14'h0ECD: rddata <= 8'hC9; 14'h0ECE: rddata <= 8'hF1; 14'h0ECF: rddata <= 8'h11;
            14'h0ED0: rddata <= 8'h1A; 14'h0ED1: rddata <= 8'h00; 14'h0ED2: rddata <= 8'hCA; 14'h0ED3: rddata <= 8'hDB;
            14'h0ED4: rddata <= 8'h03; 14'h0ED5: rddata <= 8'hBF; 14'h0ED6: rddata <= 8'hF5; 14'h0ED7: rddata <= 8'h01;
            14'h0ED8: rddata <= 8'hB5; 14'h0ED9: rddata <= 8'h0E; 14'h0EDA: rddata <= 8'hC5; 14'h0EDB: rddata <= 8'h2A;
            14'h0EDC: rddata <= 8'hAD; 14'h0EDD: rddata <= 8'h38; 14'h0EDE: rddata <= 8'h22; 14'h0EDF: rddata <= 8'hC1;
            14'h0EE0: rddata <= 8'h38; 14'h0EE1: rddata <= 8'h21; 14'h0EE2: rddata <= 8'h00; 14'h0EE3: rddata <= 8'h00;
            14'h0EE4: rddata <= 8'hE5; 14'h0EE5: rddata <= 8'h2A; 14'h0EE6: rddata <= 8'hDA; 14'h0EE7: rddata <= 8'h38;
            14'h0EE8: rddata <= 8'hE5; 14'h0EE9: rddata <= 8'h21; 14'h0EEA: rddata <= 8'hB1; 14'h0EEB: rddata <= 8'h38;
            14'h0EEC: rddata <= 8'hED; 14'h0EED: rddata <= 8'h5B; 14'h0EEE: rddata <= 8'hAF; 14'h0EEF: rddata <= 8'h38;
            14'h0EF0: rddata <= 8'hE7; 14'h0EF1: rddata <= 8'h01; 14'h0EF2: rddata <= 8'hEC; 14'h0EF3: rddata <= 8'h0E;
            14'h0EF4: rddata <= 8'hC2; 14'h0EF5: rddata <= 8'h32; 14'h0EF6: rddata <= 8'h0F; 14'h0EF7: rddata <= 8'h2A;
            14'h0EF8: rddata <= 8'hD6; 14'h0EF9: rddata <= 8'h38; 14'h0EFA: rddata <= 8'hED; 14'h0EFB: rddata <= 8'h5B;
            14'h0EFC: rddata <= 8'hD8; 14'h0EFD: rddata <= 8'h38; 14'h0EFE: rddata <= 8'hE7; 14'h0EFF: rddata <= 8'h28;
            14'h0F00: rddata <= 8'h0A; 14'h0F01: rddata <= 8'h23; 14'h0F02: rddata <= 8'h7E; 14'h0F03: rddata <= 8'h23;
            14'h0F04: rddata <= 8'hB7; 14'h0F05: rddata <= 8'hCD; 14'h0F06: rddata <= 8'h35; 14'h0F07: rddata <= 8'h0F;
            14'h0F08: rddata <= 8'h18; 14'h0F09: rddata <= 8'hF0; 14'h0F0A: rddata <= 8'hC1; 14'h0F0B: rddata <= 8'hED;
            14'h0F0C: rddata <= 8'h5B; 14'h0F0D: rddata <= 8'hDA; 14'h0F0E: rddata <= 8'h38; 14'h0F0F: rddata <= 8'hE7;
            14'h0F10: rddata <= 8'hCA; 14'h0F11: rddata <= 8'h57; 14'h0F12: rddata <= 8'h0F; 14'h0F13: rddata <= 8'hCD;
            14'h0F14: rddata <= 8'h31; 14'h0F15: rddata <= 8'h15; 14'h0F16: rddata <= 8'h7A; 14'h0F17: rddata <= 8'hE5;
            14'h0F18: rddata <= 8'h09; 14'h0F19: rddata <= 8'hB7; 14'h0F1A: rddata <= 8'hF2; 14'h0F1B: rddata <= 8'h0A;
            14'h0F1C: rddata <= 8'h0F; 14'h0F1D: rddata <= 8'h22; 14'h0F1E: rddata <= 8'hC5; 14'h0F1F: rddata <= 8'h38;
            14'h0F20: rddata <= 8'hE1; 14'h0F21: rddata <= 8'h4E; 14'h0F22: rddata <= 8'h06; 14'h0F23: rddata <= 8'h00;
            14'h0F24: rddata <= 8'h09; 14'h0F25: rddata <= 8'h09; 14'h0F26: rddata <= 8'h23; 14'h0F27: rddata <= 8'hEB;
            14'h0F28: rddata <= 8'h2A; 14'h0F29: rddata <= 8'hC5; 14'h0F2A: rddata <= 8'h38; 14'h0F2B: rddata <= 8'hEB;
            14'h0F2C: rddata <= 8'hE7; 14'h0F2D: rddata <= 8'h28; 14'h0F2E: rddata <= 8'hDC; 14'h0F2F: rddata <= 8'h01;
            14'h0F30: rddata <= 8'h27; 14'h0F31: rddata <= 8'h0F; 14'h0F32: rddata <= 8'hC5; 14'h0F33: rddata <= 8'hF6;
            14'h0F34: rddata <= 8'h80; 14'h0F35: rddata <= 8'h7E; 14'h0F36: rddata <= 8'h23; 14'h0F37: rddata <= 8'h23;
            14'h0F38: rddata <= 8'h5E; 14'h0F39: rddata <= 8'h23; 14'h0F3A: rddata <= 8'h56; 14'h0F3B: rddata <= 8'h23;
            14'h0F3C: rddata <= 8'hF0; 14'h0F3D: rddata <= 8'hB7; 14'h0F3E: rddata <= 8'hC8; 14'h0F3F: rddata <= 8'h44;
            14'h0F40: rddata <= 8'h4D; 14'h0F41: rddata <= 8'h2A; 14'h0F42: rddata <= 8'hC1; 14'h0F43: rddata <= 8'h38;
            14'h0F44: rddata <= 8'hE7; 14'h0F45: rddata <= 8'h60; 14'h0F46: rddata <= 8'h69; 14'h0F47: rddata <= 8'hD8;
            14'h0F48: rddata <= 8'hE1; 14'h0F49: rddata <= 8'hE3; 14'h0F4A: rddata <= 8'hE7; 14'h0F4B: rddata <= 8'hE3;
            14'h0F4C: rddata <= 8'hE5; 14'h0F4D: rddata <= 8'h60; 14'h0F4E: rddata <= 8'h69; 14'h0F4F: rddata <= 8'hD0;
            14'h0F50: rddata <= 8'hC1; 14'h0F51: rddata <= 8'hF1; 14'h0F52: rddata <= 8'hF1; 14'h0F53: rddata <= 8'hE5;
            14'h0F54: rddata <= 8'hD5; 14'h0F55: rddata <= 8'hC5; 14'h0F56: rddata <= 8'hC9; 14'h0F57: rddata <= 8'hD1;
            14'h0F58: rddata <= 8'hE1; 14'h0F59: rddata <= 8'h7C; 14'h0F5A: rddata <= 8'hB5; 14'h0F5B: rddata <= 8'hC8;
            14'h0F5C: rddata <= 8'h2B; 14'h0F5D: rddata <= 8'h46; 14'h0F5E: rddata <= 8'h2B; 14'h0F5F: rddata <= 8'h4E;
            14'h0F60: rddata <= 8'hE5; 14'h0F61: rddata <= 8'h2B; 14'h0F62: rddata <= 8'h2B; 14'h0F63: rddata <= 8'h6E;
            14'h0F64: rddata <= 8'h26; 14'h0F65: rddata <= 8'h00; 14'h0F66: rddata <= 8'h09; 14'h0F67: rddata <= 8'h50;
            14'h0F68: rddata <= 8'h59; 14'h0F69: rddata <= 8'h2B; 14'h0F6A: rddata <= 8'h44; 14'h0F6B: rddata <= 8'h4D;
            14'h0F6C: rddata <= 8'h2A; 14'h0F6D: rddata <= 8'hC1; 14'h0F6E: rddata <= 8'h38; 14'h0F6F: rddata <= 8'hCD;
            14'h0F70: rddata <= 8'h95; 14'h0F71: rddata <= 8'h0B; 14'h0F72: rddata <= 8'hE1; 14'h0F73: rddata <= 8'h71;
            14'h0F74: rddata <= 8'h23; 14'h0F75: rddata <= 8'h70; 14'h0F76: rddata <= 8'h60; 14'h0F77: rddata <= 8'h69;
            14'h0F78: rddata <= 8'h2B; 14'h0F79: rddata <= 8'hC3; 14'h0F7A: rddata <= 8'hDE; 14'h0F7B: rddata <= 8'h0E;
            14'h0F7C: rddata <= 8'hC5; 14'h0F7D: rddata <= 8'hE5; 14'h0F7E: rddata <= 8'h2A; 14'h0F7F: rddata <= 8'hE4;
            14'h0F80: rddata <= 8'h38; 14'h0F81: rddata <= 8'hE3; 14'h0F82: rddata <= 8'hCD; 14'h0F83: rddata <= 8'hFD;
            14'h0F84: rddata <= 8'h09; 14'h0F85: rddata <= 8'hE3; 14'h0F86: rddata <= 8'hCD; 14'h0F87: rddata <= 8'h76;
            14'h0F88: rddata <= 8'h09; 14'h0F89: rddata <= 8'h7E; 14'h0F8A: rddata <= 8'hE5; 14'h0F8B: rddata <= 8'h2A;
            14'h0F8C: rddata <= 8'hE4; 14'h0F8D: rddata <= 8'h38; 14'h0F8E: rddata <= 8'hE5; 14'h0F8F: rddata <= 8'h86;
            14'h0F90: rddata <= 8'h11; 14'h0F91: rddata <= 8'h1C; 14'h0F92: rddata <= 8'h00; 14'h0F93: rddata <= 8'hDA;
            14'h0F94: rddata <= 8'hDB; 14'h0F95: rddata <= 8'h03; 14'h0F96: rddata <= 8'hCD; 14'h0F97: rddata <= 8'h50;
            14'h0F98: rddata <= 8'h0E; 14'h0F99: rddata <= 8'hD1; 14'h0F9A: rddata <= 8'hCD; 14'h0F9B: rddata <= 8'hCD;
            14'h0F9C: rddata <= 8'h0F; 14'h0F9D: rddata <= 8'hE3; 14'h0F9E: rddata <= 8'hCD; 14'h0F9F: rddata <= 8'hCC;
            14'h0FA0: rddata <= 8'h0F; 14'h0FA1: rddata <= 8'hE5; 14'h0FA2: rddata <= 8'h2A; 14'h0FA3: rddata <= 8'hBF;
            14'h0FA4: rddata <= 8'h38; 14'h0FA5: rddata <= 8'hEB; 14'h0FA6: rddata <= 8'hCD; 14'h0FA7: rddata <= 8'hB4;
            14'h0FA8: rddata <= 8'h0F; 14'h0FA9: rddata <= 8'hCD; 14'h0FAA: rddata <= 8'hB4; 14'h0FAB: rddata <= 8'h0F;
            14'h0FAC: rddata <= 8'h21; 14'h0FAD: rddata <= 8'h91; 14'h0FAE: rddata <= 8'h09; 14'h0FAF: rddata <= 8'hE3;
            14'h0FB0: rddata <= 8'hE5; 14'h0FB1: rddata <= 8'hC3; 14'h0FB2: rddata <= 8'h7E; 14'h0FB3: rddata <= 8'h0E;
            14'h0FB4: rddata <= 8'hE1; 14'h0FB5: rddata <= 8'hE3; 14'h0FB6: rddata <= 8'h7E; 14'h0FB7: rddata <= 8'h23;
            14'h0FB8: rddata <= 8'h23; 14'h0FB9: rddata <= 8'h4E; 14'h0FBA: rddata <= 8'h23; 14'h0FBB: rddata <= 8'h46;
            14'h0FBC: rddata <= 8'h6F; 14'h0FBD: rddata <= 8'h2C; 14'h0FBE: rddata <= 8'h2D; 14'h0FBF: rddata <= 8'hC8;
            14'h0FC0: rddata <= 8'h0A; 14'h0FC1: rddata <= 8'h12; 14'h0FC2: rddata <= 8'h03; 14'h0FC3: rddata <= 8'h13;
            14'h0FC4: rddata <= 8'h18; 14'h0FC5: rddata <= 8'hF8; 14'h0FC6: rddata <= 8'hCD; 14'h0FC7: rddata <= 8'h76;
            14'h0FC8: rddata <= 8'h09; 14'h0FC9: rddata <= 8'h2A; 14'h0FCA: rddata <= 8'hE4; 14'h0FCB: rddata <= 8'h38;
            14'h0FCC: rddata <= 8'hEB; 14'h0FCD: rddata <= 8'hCD; 14'h0FCE: rddata <= 8'hE4; 14'h0FCF: rddata <= 8'h0F;
            14'h0FD0: rddata <= 8'hEB; 14'h0FD1: rddata <= 8'hC0; 14'h0FD2: rddata <= 8'hD5; 14'h0FD3: rddata <= 8'h50;
            14'h0FD4: rddata <= 8'h59; 14'h0FD5: rddata <= 8'h1B; 14'h0FD6: rddata <= 8'h4E; 14'h0FD7: rddata <= 8'h2A;
            14'h0FD8: rddata <= 8'hC1; 14'h0FD9: rddata <= 8'h38; 14'h0FDA: rddata <= 8'hE7; 14'h0FDB: rddata <= 8'h20;
            14'h0FDC: rddata <= 8'h05; 14'h0FDD: rddata <= 8'h47; 14'h0FDE: rddata <= 8'h09; 14'h0FDF: rddata <= 8'h22;
            14'h0FE0: rddata <= 8'hC1; 14'h0FE1: rddata <= 8'h38; 14'h0FE2: rddata <= 8'hE1; 14'h0FE3: rddata <= 8'hC9;
            14'h0FE4: rddata <= 8'h2A; 14'h0FE5: rddata <= 8'hAF; 14'h0FE6: rddata <= 8'h38; 14'h0FE7: rddata <= 8'h2B;
            14'h0FE8: rddata <= 8'h46; 14'h0FE9: rddata <= 8'h2B; 14'h0FEA: rddata <= 8'h4E; 14'h0FEB: rddata <= 8'h2B;
            14'h0FEC: rddata <= 8'h2B; 14'h0FED: rddata <= 8'hE7; 14'h0FEE: rddata <= 8'hC0; 14'h0FEF: rddata <= 8'h22;
            14'h0FF0: rddata <= 8'hAF; 14'h0FF1: rddata <= 8'h38; 14'h0FF2: rddata <= 8'hC9; 14'h0FF3: rddata <= 8'h01;
            14'h0FF4: rddata <= 8'h36; 14'h0FF5: rddata <= 8'h0B; 14'h0FF6: rddata <= 8'hC5; 14'h0FF7: rddata <= 8'hCD;
            14'h0FF8: rddata <= 8'hC6; 14'h0FF9: rddata <= 8'h0F; 14'h0FFA: rddata <= 8'hAF; 14'h0FFB: rddata <= 8'h57;
            14'h0FFC: rddata <= 8'h32; 14'h0FFD: rddata <= 8'hAB; 14'h0FFE: rddata <= 8'h38; 14'h0FFF: rddata <= 8'h7E;
            14'h1000: rddata <= 8'hB7; 14'h1001: rddata <= 8'hC9; 14'h1002: rddata <= 8'h01; 14'h1003: rddata <= 8'h36;
            14'h1004: rddata <= 8'h0B; 14'h1005: rddata <= 8'hC5; 14'h1006: rddata <= 8'hCD; 14'h1007: rddata <= 8'hF7;
            14'h1008: rddata <= 8'h0F; 14'h1009: rddata <= 8'hCA; 14'h100A: rddata <= 8'h97; 14'h100B: rddata <= 8'h06;
            14'h100C: rddata <= 8'h23; 14'h100D: rddata <= 8'h23; 14'h100E: rddata <= 8'h5E; 14'h100F: rddata <= 8'h23;
            14'h1010: rddata <= 8'h56; 14'h1011: rddata <= 8'h1A; 14'h1012: rddata <= 8'hC9; 14'h1013: rddata <= 8'hCD;
            14'h1014: rddata <= 8'h4E; 14'h1015: rddata <= 8'h0E; 14'h1016: rddata <= 8'hCD; 14'h1017: rddata <= 8'h57;
            14'h1018: rddata <= 8'h0B; 14'h1019: rddata <= 8'h2A; 14'h101A: rddata <= 8'hBF; 14'h101B: rddata <= 8'h38;
            14'h101C: rddata <= 8'h73; 14'h101D: rddata <= 8'hC1; 14'h101E: rddata <= 8'hC3; 14'h101F: rddata <= 8'h7E;
            14'h1020: rddata <= 8'h0E; 14'h1021: rddata <= 8'hCD; 14'h1022: rddata <= 8'hA0; 14'h1023: rddata <= 8'h10;
            14'h1024: rddata <= 8'hAF; 14'h1025: rddata <= 8'hE3; 14'h1026: rddata <= 8'h4F; 14'h1027: rddata <= 8'hE5;
            14'h1028: rddata <= 8'h7E; 14'h1029: rddata <= 8'hB8; 14'h102A: rddata <= 8'h38; 14'h102B: rddata <= 8'h02;
            14'h102C: rddata <= 8'h78; 14'h102D: rddata <= 8'h11; 14'h102E: rddata <= 8'h0E; 14'h102F: rddata <= 8'h00;
            14'h1030: rddata <= 8'hC5; 14'h1031: rddata <= 8'hCD; 14'h1032: rddata <= 8'hB3; 14'h1033: rddata <= 8'h0E;
            14'h1034: rddata <= 8'hC1; 14'h1035: rddata <= 8'hE1; 14'h1036: rddata <= 8'hE5; 14'h1037: rddata <= 8'h23;
            14'h1038: rddata <= 8'h23; 14'h1039: rddata <= 8'h46; 14'h103A: rddata <= 8'h23; 14'h103B: rddata <= 8'h66;
            14'h103C: rddata <= 8'h68; 14'h103D: rddata <= 8'h06; 14'h103E: rddata <= 8'h00; 14'h103F: rddata <= 8'h09;
            14'h1040: rddata <= 8'h44; 14'h1041: rddata <= 8'h4D; 14'h1042: rddata <= 8'hCD; 14'h1043: rddata <= 8'h53;
            14'h1044: rddata <= 8'h0E; 14'h1045: rddata <= 8'h6F; 14'h1046: rddata <= 8'hCD; 14'h1047: rddata <= 8'hBD;
            14'h1048: rddata <= 8'h0F; 14'h1049: rddata <= 8'hD1; 14'h104A: rddata <= 8'hCD; 14'h104B: rddata <= 8'hCD;
            14'h104C: rddata <= 8'h0F; 14'h104D: rddata <= 8'hC3; 14'h104E: rddata <= 8'h7E; 14'h104F: rddata <= 8'h0E;
            14'h1050: rddata <= 8'hCD; 14'h1051: rddata <= 8'hA0; 14'h1052: rddata <= 8'h10; 14'h1053: rddata <= 8'hD1;
            14'h1054: rddata <= 8'hD5; 14'h1055: rddata <= 8'h1A; 14'h1056: rddata <= 8'h90; 14'h1057: rddata <= 8'h18;
            14'h1058: rddata <= 8'hCC; 14'h1059: rddata <= 8'hEB; 14'h105A: rddata <= 8'h7E; 14'h105B: rddata <= 8'hCD;
            14'h105C: rddata <= 8'hA3; 14'h105D: rddata <= 8'h10; 14'h105E: rddata <= 8'h04; 14'h105F: rddata <= 8'h05;
            14'h1060: rddata <= 8'hCA; 14'h1061: rddata <= 8'h97; 14'h1062: rddata <= 8'h06; 14'h1063: rddata <= 8'hC5;
            14'h1064: rddata <= 8'h1E; 14'h1065: rddata <= 8'hFF; 14'h1066: rddata <= 8'hFE; 14'h1067: rddata <= 8'h29;
            14'h1068: rddata <= 8'h28; 14'h1069: rddata <= 8'h05; 14'h106A: rddata <= 8'hCF; 14'h106B: rddata <= 8'h2C;
            14'h106C: rddata <= 8'hCD; 14'h106D: rddata <= 8'h54; 14'h106E: rddata <= 8'h0B; 14'h106F: rddata <= 8'hCF;
            14'h1070: rddata <= 8'h29; 14'h1071: rddata <= 8'hF1; 14'h1072: rddata <= 8'hE3; 14'h1073: rddata <= 8'h01;
            14'h1074: rddata <= 8'h27; 14'h1075: rddata <= 8'h10; 14'h1076: rddata <= 8'hC5; 14'h1077: rddata <= 8'h3D;
            14'h1078: rddata <= 8'hBE; 14'h1079: rddata <= 8'h06; 14'h107A: rddata <= 8'h00; 14'h107B: rddata <= 8'hD0;
            14'h107C: rddata <= 8'h4F; 14'h107D: rddata <= 8'h7E; 14'h107E: rddata <= 8'h91; 14'h107F: rddata <= 8'hBB;
            14'h1080: rddata <= 8'h47; 14'h1081: rddata <= 8'hD8; 14'h1082: rddata <= 8'h43; 14'h1083: rddata <= 8'hC9;
            14'h1084: rddata <= 8'hCD; 14'h1085: rddata <= 8'hF7; 14'h1086: rddata <= 8'h0F; 14'h1087: rddata <= 8'hCA;
            14'h1088: rddata <= 8'hC3; 14'h1089: rddata <= 8'h12; 14'h108A: rddata <= 8'h5F; 14'h108B: rddata <= 8'h23;
            14'h108C: rddata <= 8'h23; 14'h108D: rddata <= 8'h7E; 14'h108E: rddata <= 8'h23; 14'h108F: rddata <= 8'h66;
            14'h1090: rddata <= 8'h6F; 14'h1091: rddata <= 8'hE5; 14'h1092: rddata <= 8'h19; 14'h1093: rddata <= 8'h46;
            14'h1094: rddata <= 8'h72; 14'h1095: rddata <= 8'hE3; 14'h1096: rddata <= 8'hC5; 14'h1097: rddata <= 8'h2B;
            14'h1098: rddata <= 8'hD7; 14'h1099: rddata <= 8'hCD; 14'h109A: rddata <= 8'hE5; 14'h109B: rddata <= 8'h15;
            14'h109C: rddata <= 8'hC1; 14'h109D: rddata <= 8'hE1; 14'h109E: rddata <= 8'h70; 14'h109F: rddata <= 8'hC9;
            14'h10A0: rddata <= 8'hEB; 14'h10A1: rddata <= 8'hCF; 14'h10A2: rddata <= 8'h29; 14'h10A3: rddata <= 8'hC1;
            14'h10A4: rddata <= 8'hD1; 14'h10A5: rddata <= 8'hC5; 14'h10A6: rddata <= 8'h43; 14'h10A7: rddata <= 8'hC9;
            14'h10A8: rddata <= 8'h2A; 14'h10A9: rddata <= 8'hDA; 14'h10AA: rddata <= 8'h38; 14'h10AB: rddata <= 8'hEB;
            14'h10AC: rddata <= 8'h21; 14'h10AD: rddata <= 8'h00; 14'h10AE: rddata <= 8'h00; 14'h10AF: rddata <= 8'h39;
            14'h10B0: rddata <= 8'h3A; 14'h10B1: rddata <= 8'hAB; 14'h10B2: rddata <= 8'h38; 14'h10B3: rddata <= 8'hB7;
            14'h10B4: rddata <= 8'hCA; 14'h10B5: rddata <= 8'h1C; 14'h10B6: rddata <= 8'h0B; 14'h10B7: rddata <= 8'hCD;
            14'h10B8: rddata <= 8'hC9; 14'h10B9: rddata <= 8'h0F; 14'h10BA: rddata <= 8'hCD; 14'h10BB: rddata <= 8'hDB;
            14'h10BC: rddata <= 8'h0E; 14'h10BD: rddata <= 8'hED; 14'h10BE: rddata <= 8'h5B; 14'h10BF: rddata <= 8'h4B;
            14'h10C0: rddata <= 8'h38; 14'h10C1: rddata <= 8'h2A; 14'h10C2: rddata <= 8'hC1; 14'h10C3: rddata <= 8'h38;
            14'h10C4: rddata <= 8'hC3; 14'h10C5: rddata <= 8'h1C; 14'h10C6: rddata <= 8'h0B; 14'h10C7: rddata <= 8'h2B;
            14'h10C8: rddata <= 8'hD7; 14'h10C9: rddata <= 8'hC8; 14'h10CA: rddata <= 8'hCF; 14'h10CB: rddata <= 8'h2C;
            14'h10CC: rddata <= 8'h01; 14'h10CD: rddata <= 8'hC7; 14'h10CE: rddata <= 8'h10; 14'h10CF: rddata <= 8'hC5;
            14'h10D0: rddata <= 8'hF6; 14'h10D1: rddata <= 8'hAF; 14'h10D2: rddata <= 8'h32; 14'h10D3: rddata <= 8'hAA;
            14'h10D4: rddata <= 8'h38; 14'h10D5: rddata <= 8'h4E; 14'h10D6: rddata <= 8'hCD; 14'h10D7: rddata <= 8'hC5;
            14'h10D8: rddata <= 8'h0C; 14'h10D9: rddata <= 8'hDA; 14'h10DA: rddata <= 8'hC4; 14'h10DB: rddata <= 8'h03;
            14'h10DC: rddata <= 8'hAF; 14'h10DD: rddata <= 8'h47; 14'h10DE: rddata <= 8'h32; 14'h10DF: rddata <= 8'hAB;
            14'h10E0: rddata <= 8'h38; 14'h10E1: rddata <= 8'hD7; 14'h10E2: rddata <= 8'h38; 14'h10E3: rddata <= 8'h05;
            14'h10E4: rddata <= 8'hCD; 14'h10E5: rddata <= 8'hC6; 14'h10E6: rddata <= 8'h0C; 14'h10E7: rddata <= 8'h38;
            14'h10E8: rddata <= 8'h09; 14'h10E9: rddata <= 8'h47; 14'h10EA: rddata <= 8'hD7; 14'h10EB: rddata <= 8'h38;
            14'h10EC: rddata <= 8'hFD; 14'h10ED: rddata <= 8'hCD; 14'h10EE: rddata <= 8'hC6; 14'h10EF: rddata <= 8'h0C;
            14'h10F0: rddata <= 8'h30; 14'h10F1: rddata <= 8'hF8; 14'h10F2: rddata <= 8'hD6; 14'h10F3: rddata <= 8'h24;
            14'h10F4: rddata <= 8'h20; 14'h10F5: rddata <= 8'h08; 14'h10F6: rddata <= 8'h3C; 14'h10F7: rddata <= 8'h32;
            14'h10F8: rddata <= 8'hAB; 14'h10F9: rddata <= 8'h38; 14'h10FA: rddata <= 8'h0F; 14'h10FB: rddata <= 8'h80;
            14'h10FC: rddata <= 8'h47; 14'h10FD: rddata <= 8'hD7; 14'h10FE: rddata <= 8'h3A; 14'h10FF: rddata <= 8'hCB;
            14'h1100: rddata <= 8'h38; 14'h1101: rddata <= 8'h3D; 14'h1102: rddata <= 8'hCA; 14'h1103: rddata <= 8'hA0;
            14'h1104: rddata <= 8'h11; 14'h1105: rddata <= 8'hF2; 14'h1106: rddata <= 8'h0E; 14'h1107: rddata <= 8'h11;
            14'h1108: rddata <= 8'h7E; 14'h1109: rddata <= 8'hD6; 14'h110A: rddata <= 8'h28; 14'h110B: rddata <= 8'hCA;
            14'h110C: rddata <= 8'h7A; 14'h110D: rddata <= 8'h11; 14'h110E: rddata <= 8'hAF; 14'h110F: rddata <= 8'h32;
            14'h1110: rddata <= 8'hCB; 14'h1111: rddata <= 8'h38; 14'h1112: rddata <= 8'hE5; 14'h1113: rddata <= 8'h50;
            14'h1114: rddata <= 8'h59; 14'h1115: rddata <= 8'h2A; 14'h1116: rddata <= 8'hDE; 14'h1117: rddata <= 8'h38;
            14'h1118: rddata <= 8'hE7; 14'h1119: rddata <= 8'h11; 14'h111A: rddata <= 8'hE0; 14'h111B: rddata <= 8'h38;
            14'h111C: rddata <= 8'hCA; 14'h111D: rddata <= 8'h1A; 14'h111E: rddata <= 8'h14; 14'h111F: rddata <= 8'h2A;
            14'h1120: rddata <= 8'hD8; 14'h1121: rddata <= 8'h38; 14'h1122: rddata <= 8'hEB; 14'h1123: rddata <= 8'h2A;
            14'h1124: rddata <= 8'hD6; 14'h1125: rddata <= 8'h38; 14'h1126: rddata <= 8'hE7; 14'h1127: rddata <= 8'hCA;
            14'h1128: rddata <= 8'h3D; 14'h1129: rddata <= 8'h11; 14'h112A: rddata <= 8'h79; 14'h112B: rddata <= 8'h96;
            14'h112C: rddata <= 8'h23; 14'h112D: rddata <= 8'hC2; 14'h112E: rddata <= 8'h32; 14'h112F: rddata <= 8'h11;
            14'h1130: rddata <= 8'h78; 14'h1131: rddata <= 8'h96; 14'h1132: rddata <= 8'h23; 14'h1133: rddata <= 8'hCA;
            14'h1134: rddata <= 8'h6C; 14'h1135: rddata <= 8'h11; 14'h1136: rddata <= 8'h23; 14'h1137: rddata <= 8'h23;
            14'h1138: rddata <= 8'h23; 14'h1139: rddata <= 8'h23; 14'h113A: rddata <= 8'hC3; 14'h113B: rddata <= 8'h26;
            14'h113C: rddata <= 8'h11; 14'h113D: rddata <= 8'hE1; 14'h113E: rddata <= 8'hE3; 14'h113F: rddata <= 8'hD5;
            14'h1140: rddata <= 8'h11; 14'h1141: rddata <= 8'h51; 14'h1142: rddata <= 8'h0A; 14'h1143: rddata <= 8'hE7;
            14'h1144: rddata <= 8'hD1; 14'h1145: rddata <= 8'hCA; 14'h1146: rddata <= 8'h6F; 14'h1147: rddata <= 8'h11;
            14'h1148: rddata <= 8'hE3; 14'h1149: rddata <= 8'hE5; 14'h114A: rddata <= 8'hC5; 14'h114B: rddata <= 8'h01;
            14'h114C: rddata <= 8'h06; 14'h114D: rddata <= 8'h00; 14'h114E: rddata <= 8'h2A; 14'h114F: rddata <= 8'hDA;
            14'h1150: rddata <= 8'h38; 14'h1151: rddata <= 8'hE5; 14'h1152: rddata <= 8'h09; 14'h1153: rddata <= 8'hC1;
            14'h1154: rddata <= 8'hE5; 14'h1155: rddata <= 8'hCD; 14'h1156: rddata <= 8'h92; 14'h1157: rddata <= 8'h0B;
            14'h1158: rddata <= 8'hE1; 14'h1159: rddata <= 8'h22; 14'h115A: rddata <= 8'hDA; 14'h115B: rddata <= 8'h38;
            14'h115C: rddata <= 8'h60; 14'h115D: rddata <= 8'h69; 14'h115E: rddata <= 8'h22; 14'h115F: rddata <= 8'hD8;
            14'h1160: rddata <= 8'h38; 14'h1161: rddata <= 8'h2B; 14'h1162: rddata <= 8'h36; 14'h1163: rddata <= 8'h00;
            14'h1164: rddata <= 8'hE7; 14'h1165: rddata <= 8'h20; 14'h1166: rddata <= 8'hFA; 14'h1167: rddata <= 8'hD1;
            14'h1168: rddata <= 8'h73; 14'h1169: rddata <= 8'h23; 14'h116A: rddata <= 8'h72; 14'h116B: rddata <= 8'h23;
            14'h116C: rddata <= 8'hEB; 14'h116D: rddata <= 8'hE1; 14'h116E: rddata <= 8'hC9; 14'h116F: rddata <= 8'h32;
            14'h1170: rddata <= 8'hE7; 14'h1171: rddata <= 8'h38; 14'h1172: rddata <= 8'h21; 14'h1173: rddata <= 8'h6D;
            14'h1174: rddata <= 8'h03; 14'h1175: rddata <= 8'h22; 14'h1176: rddata <= 8'hE4; 14'h1177: rddata <= 8'h38;
            14'h1178: rddata <= 8'hE1; 14'h1179: rddata <= 8'hC9; 14'h117A: rddata <= 8'hE5; 14'h117B: rddata <= 8'h2A;
            14'h117C: rddata <= 8'hAA; 14'h117D: rddata <= 8'h38; 14'h117E: rddata <= 8'hE3; 14'h117F: rddata <= 8'h57;
            14'h1180: rddata <= 8'hD5; 14'h1181: rddata <= 8'hC5; 14'h1182: rddata <= 8'hCD; 14'h1183: rddata <= 8'h7A;
            14'h1184: rddata <= 8'h06; 14'h1185: rddata <= 8'hC1; 14'h1186: rddata <= 8'hF1; 14'h1187: rddata <= 8'hEB;
            14'h1188: rddata <= 8'hE3; 14'h1189: rddata <= 8'hE5; 14'h118A: rddata <= 8'hEB; 14'h118B: rddata <= 8'h3C;
            14'h118C: rddata <= 8'h57; 14'h118D: rddata <= 8'h7E; 14'h118E: rddata <= 8'hFE; 14'h118F: rddata <= 8'h2C;
            14'h1190: rddata <= 8'hCA; 14'h1191: rddata <= 8'h80; 14'h1192: rddata <= 8'h11; 14'h1193: rddata <= 8'hCF;
            14'h1194: rddata <= 8'h29; 14'h1195: rddata <= 8'h22; 14'h1196: rddata <= 8'hD0; 14'h1197: rddata <= 8'h38;
            14'h1198: rddata <= 8'hE1; 14'h1199: rddata <= 8'h22; 14'h119A: rddata <= 8'hAA; 14'h119B: rddata <= 8'h38;
            14'h119C: rddata <= 8'h1E; 14'h119D: rddata <= 8'h00; 14'h119E: rddata <= 8'hD5; 14'h119F: rddata <= 8'h11;
            14'h11A0: rddata <= 8'hE5; 14'h11A1: rddata <= 8'hF5; 14'h11A2: rddata <= 8'h2A; 14'h11A3: rddata <= 8'hD8;
            14'h11A4: rddata <= 8'h38; 14'h11A5: rddata <= 8'h3E; 14'h11A6: rddata <= 8'h19; 14'h11A7: rddata <= 8'hED;
            14'h11A8: rddata <= 8'h5B; 14'h11A9: rddata <= 8'hDA; 14'h11AA: rddata <= 8'h38; 14'h11AB: rddata <= 8'hE7;
            14'h11AC: rddata <= 8'h28; 14'h11AD: rddata <= 8'h25; 14'h11AE: rddata <= 8'h7E; 14'h11AF: rddata <= 8'h23;
            14'h11B0: rddata <= 8'hB9; 14'h11B1: rddata <= 8'h20; 14'h11B2: rddata <= 8'h02; 14'h11B3: rddata <= 8'h7E;
            14'h11B4: rddata <= 8'hB8; 14'h11B5: rddata <= 8'h23; 14'h11B6: rddata <= 8'h5E; 14'h11B7: rddata <= 8'h23;
            14'h11B8: rddata <= 8'h56; 14'h11B9: rddata <= 8'h23; 14'h11BA: rddata <= 8'h20; 14'h11BB: rddata <= 8'hEA;
            14'h11BC: rddata <= 8'h3A; 14'h11BD: rddata <= 8'hAA; 14'h11BE: rddata <= 8'h38; 14'h11BF: rddata <= 8'hB7;
            14'h11C0: rddata <= 8'hC2; 14'h11C1: rddata <= 8'hCD; 14'h11C2: rddata <= 8'h03; 14'h11C3: rddata <= 8'hF1;
            14'h11C4: rddata <= 8'h44; 14'h11C5: rddata <= 8'h4D; 14'h11C6: rddata <= 8'hCA; 14'h11C7: rddata <= 8'h1A;
            14'h11C8: rddata <= 8'h14; 14'h11C9: rddata <= 8'h96; 14'h11CA: rddata <= 8'hCA; 14'h11CB: rddata <= 8'h2B;
            14'h11CC: rddata <= 8'h12; 14'h11CD: rddata <= 8'h11; 14'h11CE: rddata <= 8'h10; 14'h11CF: rddata <= 8'h00;
            14'h11D0: rddata <= 8'hC3; 14'h11D1: rddata <= 8'hDB; 14'h11D2: rddata <= 8'h03; 14'h11D3: rddata <= 8'h11;
            14'h11D4: rddata <= 8'h04; 14'h11D5: rddata <= 8'h00; 14'h11D6: rddata <= 8'hF1; 14'h11D7: rddata <= 8'hCA;
            14'h11D8: rddata <= 8'h97; 14'h11D9: rddata <= 8'h06; 14'h11DA: rddata <= 8'h71; 14'h11DB: rddata <= 8'h23;
            14'h11DC: rddata <= 8'h70; 14'h11DD: rddata <= 8'h23; 14'h11DE: rddata <= 8'h4F; 14'h11DF: rddata <= 8'hCD;
            14'h11E0: rddata <= 8'hA0; 14'h11E1: rddata <= 8'h0B; 14'h11E2: rddata <= 8'h23; 14'h11E3: rddata <= 8'h23;
            14'h11E4: rddata <= 8'h22; 14'h11E5: rddata <= 8'hC3; 14'h11E6: rddata <= 8'h38; 14'h11E7: rddata <= 8'h71;
            14'h11E8: rddata <= 8'h23; 14'h11E9: rddata <= 8'h3A; 14'h11EA: rddata <= 8'hAA; 14'h11EB: rddata <= 8'h38;
            14'h11EC: rddata <= 8'h17; 14'h11ED: rddata <= 8'h79; 14'h11EE: rddata <= 8'h01; 14'h11EF: rddata <= 8'h0B;
            14'h11F0: rddata <= 8'h00; 14'h11F1: rddata <= 8'h30; 14'h11F2: rddata <= 8'h02; 14'h11F3: rddata <= 8'hC1;
            14'h11F4: rddata <= 8'h03; 14'h11F5: rddata <= 8'h71; 14'h11F6: rddata <= 8'hF5; 14'h11F7: rddata <= 8'h23;
            14'h11F8: rddata <= 8'h70; 14'h11F9: rddata <= 8'h23; 14'h11FA: rddata <= 8'hE5; 14'h11FB: rddata <= 8'hCD;
            14'h11FC: rddata <= 8'hCA; 14'h11FD: rddata <= 8'h15; 14'h11FE: rddata <= 8'hEB; 14'h11FF: rddata <= 8'hE1;
            14'h1200: rddata <= 8'hF1; 14'h1201: rddata <= 8'h3D; 14'h1202: rddata <= 8'h20; 14'h1203: rddata <= 8'hEA;
            14'h1204: rddata <= 8'hF5; 14'h1205: rddata <= 8'h42; 14'h1206: rddata <= 8'h4B; 14'h1207: rddata <= 8'hEB;
            14'h1208: rddata <= 8'h19; 14'h1209: rddata <= 8'hDA; 14'h120A: rddata <= 8'hB7; 14'h120B: rddata <= 8'h0B;
            14'h120C: rddata <= 8'hCD; 14'h120D: rddata <= 8'hA9; 14'h120E: rddata <= 8'h0B; 14'h120F: rddata <= 8'h22;
            14'h1210: rddata <= 8'hDA; 14'h1211: rddata <= 8'h38; 14'h1212: rddata <= 8'h2B; 14'h1213: rddata <= 8'h36;
            14'h1214: rddata <= 8'h00; 14'h1215: rddata <= 8'hE7; 14'h1216: rddata <= 8'h20; 14'h1217: rddata <= 8'hFA;
            14'h1218: rddata <= 8'h03; 14'h1219: rddata <= 8'h57; 14'h121A: rddata <= 8'h2A; 14'h121B: rddata <= 8'hC3;
            14'h121C: rddata <= 8'h38; 14'h121D: rddata <= 8'h5E; 14'h121E: rddata <= 8'hEB; 14'h121F: rddata <= 8'h29;
            14'h1220: rddata <= 8'h09; 14'h1221: rddata <= 8'hEB; 14'h1222: rddata <= 8'h2B; 14'h1223: rddata <= 8'h2B;
            14'h1224: rddata <= 8'h73; 14'h1225: rddata <= 8'h23; 14'h1226: rddata <= 8'h72; 14'h1227: rddata <= 8'h23;
            14'h1228: rddata <= 8'hF1; 14'h1229: rddata <= 8'h38; 14'h122A: rddata <= 8'h21; 14'h122B: rddata <= 8'h47;
            14'h122C: rddata <= 8'h4F; 14'h122D: rddata <= 8'h7E; 14'h122E: rddata <= 8'h23; 14'h122F: rddata <= 8'h16;
            14'h1230: rddata <= 8'hE1; 14'h1231: rddata <= 8'h5E; 14'h1232: rddata <= 8'h23; 14'h1233: rddata <= 8'h56;
            14'h1234: rddata <= 8'h23; 14'h1235: rddata <= 8'hE3; 14'h1236: rddata <= 8'hF5; 14'h1237: rddata <= 8'hE7;
            14'h1238: rddata <= 8'hD2; 14'h1239: rddata <= 8'hCD; 14'h123A: rddata <= 8'h11; 14'h123B: rddata <= 8'hE5;
            14'h123C: rddata <= 8'hCD; 14'h123D: rddata <= 8'hCA; 14'h123E: rddata <= 8'h15; 14'h123F: rddata <= 8'hD1;
            14'h1240: rddata <= 8'h19; 14'h1241: rddata <= 8'hF1; 14'h1242: rddata <= 8'h3D; 14'h1243: rddata <= 8'h44;
            14'h1244: rddata <= 8'h4D; 14'h1245: rddata <= 8'h20; 14'h1246: rddata <= 8'hE9; 14'h1247: rddata <= 8'h29;
            14'h1248: rddata <= 8'h29; 14'h1249: rddata <= 8'hC1; 14'h124A: rddata <= 8'h09; 14'h124B: rddata <= 8'hEB;
            14'h124C: rddata <= 8'h2A; 14'h124D: rddata <= 8'hD0; 14'h124E: rddata <= 8'h38; 14'h124F: rddata <= 8'hC9;
            14'h1250: rddata <= 8'h21; 14'h1251: rddata <= 8'h57; 14'h1252: rddata <= 8'h17; 14'h1253: rddata <= 8'hCD;
            14'h1254: rddata <= 8'h31; 14'h1255: rddata <= 8'h15; 14'h1256: rddata <= 8'h18; 14'h1257: rddata <= 8'h09;
            14'h1258: rddata <= 8'hCD; 14'h1259: rddata <= 8'h31; 14'h125A: rddata <= 8'h15; 14'h125B: rddata <= 8'h21;
            14'h125C: rddata <= 8'hC1; 14'h125D: rddata <= 8'hD1; 14'h125E: rddata <= 8'hCD; 14'h125F: rddata <= 8'h0B;
            14'h1260: rddata <= 8'h15; 14'h1261: rddata <= 8'h78; 14'h1262: rddata <= 8'hB7; 14'h1263: rddata <= 8'hC8;
            14'h1264: rddata <= 8'h3A; 14'h1265: rddata <= 8'hE7; 14'h1266: rddata <= 8'h38; 14'h1267: rddata <= 8'hB7;
            14'h1268: rddata <= 8'hCA; 14'h1269: rddata <= 8'h23; 14'h126A: rddata <= 8'h15; 14'h126B: rddata <= 8'h90;
            14'h126C: rddata <= 8'h30; 14'h126D: rddata <= 8'h0C; 14'h126E: rddata <= 8'h2F; 14'h126F: rddata <= 8'h3C;
            14'h1270: rddata <= 8'hEB; 14'h1271: rddata <= 8'hCD; 14'h1272: rddata <= 8'h13; 14'h1273: rddata <= 8'h15;
            14'h1274: rddata <= 8'hEB; 14'h1275: rddata <= 8'hCD; 14'h1276: rddata <= 8'h23; 14'h1277: rddata <= 8'h15;
            14'h1278: rddata <= 8'hC1; 14'h1279: rddata <= 8'hD1; 14'h127A: rddata <= 8'hFE; 14'h127B: rddata <= 8'h19;
            14'h127C: rddata <= 8'hD0; 14'h127D: rddata <= 8'hF5; 14'h127E: rddata <= 8'hCD; 14'h127F: rddata <= 8'h46;
            14'h1280: rddata <= 8'h15; 14'h1281: rddata <= 8'h67; 14'h1282: rddata <= 8'hF1; 14'h1283: rddata <= 8'hCD;
            14'h1284: rddata <= 8'h30; 14'h1285: rddata <= 8'h13; 14'h1286: rddata <= 8'h7C; 14'h1287: rddata <= 8'hB7;
            14'h1288: rddata <= 8'h21; 14'h1289: rddata <= 8'hE4; 14'h128A: rddata <= 8'h38; 14'h128B: rddata <= 8'hF2;
            14'h128C: rddata <= 8'h9F; 14'h128D: rddata <= 8'h12; 14'h128E: rddata <= 8'hCD; 14'h128F: rddata <= 8'h10;
            14'h1290: rddata <= 8'h13; 14'h1291: rddata <= 8'h30; 14'h1292: rddata <= 8'h5E; 14'h1293: rddata <= 8'h23;
            14'h1294: rddata <= 8'h34; 14'h1295: rddata <= 8'hCA; 14'h1296: rddata <= 8'hD3; 14'h1297: rddata <= 8'h03;
            14'h1298: rddata <= 8'h2E; 14'h1299: rddata <= 8'h01; 14'h129A: rddata <= 8'hCD; 14'h129B: rddata <= 8'h52;
            14'h129C: rddata <= 8'h13; 14'h129D: rddata <= 8'h18; 14'h129E: rddata <= 8'h52; 14'h129F: rddata <= 8'hAF;
            14'h12A0: rddata <= 8'h90; 14'h12A1: rddata <= 8'h47; 14'h12A2: rddata <= 8'h7E; 14'h12A3: rddata <= 8'h9B;
            14'h12A4: rddata <= 8'h5F; 14'h12A5: rddata <= 8'h23; 14'h12A6: rddata <= 8'h7E; 14'h12A7: rddata <= 8'h9A;
            14'h12A8: rddata <= 8'h57; 14'h12A9: rddata <= 8'h23; 14'h12AA: rddata <= 8'h7E; 14'h12AB: rddata <= 8'h99;
            14'h12AC: rddata <= 8'h4F; 14'h12AD: rddata <= 8'hDC; 14'h12AE: rddata <= 8'h1C; 14'h12AF: rddata <= 8'h13;
            14'h12B0: rddata <= 8'h68; 14'h12B1: rddata <= 8'h63; 14'h12B2: rddata <= 8'hAF; 14'h12B3: rddata <= 8'h47;
            14'h12B4: rddata <= 8'h79; 14'h12B5: rddata <= 8'hB7; 14'h12B6: rddata <= 8'h20; 14'h12B7: rddata <= 8'h27;
            14'h12B8: rddata <= 8'h4A; 14'h12B9: rddata <= 8'h54; 14'h12BA: rddata <= 8'h65; 14'h12BB: rddata <= 8'h6F;
            14'h12BC: rddata <= 8'h78; 14'h12BD: rddata <= 8'hD6; 14'h12BE: rddata <= 8'h08; 14'h12BF: rddata <= 8'hFE;
            14'h12C0: rddata <= 8'hE0; 14'h12C1: rddata <= 8'h20; 14'h12C2: rddata <= 8'hF0; 14'h12C3: rddata <= 8'hAF;
            14'h12C4: rddata <= 8'h32; 14'h12C5: rddata <= 8'hE7; 14'h12C6: rddata <= 8'h38; 14'h12C7: rddata <= 8'hC9;
            14'h12C8: rddata <= 8'h7C; 14'h12C9: rddata <= 8'hB5; 14'h12CA: rddata <= 8'hB2; 14'h12CB: rddata <= 8'h20;
            14'h12CC: rddata <= 8'h0A; 14'h12CD: rddata <= 8'h79; 14'h12CE: rddata <= 8'h05; 14'h12CF: rddata <= 8'h17;
            14'h12D0: rddata <= 8'h30; 14'h12D1: rddata <= 8'hFC; 14'h12D2: rddata <= 8'h04; 14'h12D3: rddata <= 8'h1F;
            14'h12D4: rddata <= 8'h4F; 14'h12D5: rddata <= 8'h18; 14'h12D6: rddata <= 8'h0B; 14'h12D7: rddata <= 8'h05;
            14'h12D8: rddata <= 8'h29; 14'h12D9: rddata <= 8'h7A; 14'h12DA: rddata <= 8'h17; 14'h12DB: rddata <= 8'h57;
            14'h12DC: rddata <= 8'h79; 14'h12DD: rddata <= 8'h8F; 14'h12DE: rddata <= 8'h4F; 14'h12DF: rddata <= 8'hF2;
            14'h12E0: rddata <= 8'hC8; 14'h12E1: rddata <= 8'h12; 14'h12E2: rddata <= 8'h78; 14'h12E3: rddata <= 8'h5C;
            14'h12E4: rddata <= 8'h45; 14'h12E5: rddata <= 8'hB7; 14'h12E6: rddata <= 8'h28; 14'h12E7: rddata <= 8'h09;
            14'h12E8: rddata <= 8'h21; 14'h12E9: rddata <= 8'hE7; 14'h12EA: rddata <= 8'h38; 14'h12EB: rddata <= 8'h86;
            14'h12EC: rddata <= 8'h77; 14'h12ED: rddata <= 8'h30; 14'h12EE: rddata <= 8'hD4; 14'h12EF: rddata <= 8'h28;
            14'h12F0: rddata <= 8'hD2; 14'h12F1: rddata <= 8'h78; 14'h12F2: rddata <= 8'h21; 14'h12F3: rddata <= 8'hE7;
            14'h12F4: rddata <= 8'h38; 14'h12F5: rddata <= 8'hB7; 14'h12F6: rddata <= 8'hFC; 14'h12F7: rddata <= 8'h03;
            14'h12F8: rddata <= 8'h13; 14'h12F9: rddata <= 8'h46; 14'h12FA: rddata <= 8'h23; 14'h12FB: rddata <= 8'h7E;
            14'h12FC: rddata <= 8'hE6; 14'h12FD: rddata <= 8'h80; 14'h12FE: rddata <= 8'hA9; 14'h12FF: rddata <= 8'h4F;
            14'h1300: rddata <= 8'hC3; 14'h1301: rddata <= 8'h23; 14'h1302: rddata <= 8'h15; 14'h1303: rddata <= 8'h1C;
            14'h1304: rddata <= 8'hC0; 14'h1305: rddata <= 8'h14; 14'h1306: rddata <= 8'hC0; 14'h1307: rddata <= 8'h0C;
            14'h1308: rddata <= 8'hC0; 14'h1309: rddata <= 8'h0E; 14'h130A: rddata <= 8'h80; 14'h130B: rddata <= 8'h34;
            14'h130C: rddata <= 8'hC0; 14'h130D: rddata <= 8'hC3; 14'h130E: rddata <= 8'hD3; 14'h130F: rddata <= 8'h03;
            14'h1310: rddata <= 8'h7E; 14'h1311: rddata <= 8'h83; 14'h1312: rddata <= 8'h5F; 14'h1313: rddata <= 8'h23;
            14'h1314: rddata <= 8'h7E; 14'h1315: rddata <= 8'h8A; 14'h1316: rddata <= 8'h57; 14'h1317: rddata <= 8'h23;
            14'h1318: rddata <= 8'h7E; 14'h1319: rddata <= 8'h89; 14'h131A: rddata <= 8'h4F; 14'h131B: rddata <= 8'hC9;
            14'h131C: rddata <= 8'h21; 14'h131D: rddata <= 8'hE8; 14'h131E: rddata <= 8'h38; 14'h131F: rddata <= 8'h7E;
            14'h1320: rddata <= 8'h2F; 14'h1321: rddata <= 8'h77; 14'h1322: rddata <= 8'hAF; 14'h1323: rddata <= 8'h6F;
            14'h1324: rddata <= 8'h90; 14'h1325: rddata <= 8'h47; 14'h1326: rddata <= 8'h7D; 14'h1327: rddata <= 8'h9B;
            14'h1328: rddata <= 8'h5F; 14'h1329: rddata <= 8'h7D; 14'h132A: rddata <= 8'h9A; 14'h132B: rddata <= 8'h57;
            14'h132C: rddata <= 8'h7D; 14'h132D: rddata <= 8'h99; 14'h132E: rddata <= 8'h4F; 14'h132F: rddata <= 8'hC9;
            14'h1330: rddata <= 8'h06; 14'h1331: rddata <= 8'h00; 14'h1332: rddata <= 8'hD6; 14'h1333: rddata <= 8'h08;
            14'h1334: rddata <= 8'h38; 14'h1335: rddata <= 8'h07; 14'h1336: rddata <= 8'h43; 14'h1337: rddata <= 8'h5A;
            14'h1338: rddata <= 8'h51; 14'h1339: rddata <= 8'h0E; 14'h133A: rddata <= 8'h00; 14'h133B: rddata <= 8'h18;
            14'h133C: rddata <= 8'hF5; 14'h133D: rddata <= 8'hC6; 14'h133E: rddata <= 8'h09; 14'h133F: rddata <= 8'h6F;
            14'h1340: rddata <= 8'h7A; 14'h1341: rddata <= 8'hB3; 14'h1342: rddata <= 8'hB0; 14'h1343: rddata <= 8'h20;
            14'h1344: rddata <= 8'h09; 14'h1345: rddata <= 8'h79; 14'h1346: rddata <= 8'h2D; 14'h1347: rddata <= 8'hC8;
            14'h1348: rddata <= 8'h1F; 14'h1349: rddata <= 8'h4F; 14'h134A: rddata <= 8'h30; 14'h134B: rddata <= 8'hFA;
            14'h134C: rddata <= 8'h18; 14'h134D: rddata <= 8'h06; 14'h134E: rddata <= 8'hAF; 14'h134F: rddata <= 8'h2D;
            14'h1350: rddata <= 8'hC8; 14'h1351: rddata <= 8'h79; 14'h1352: rddata <= 8'h1F; 14'h1353: rddata <= 8'h4F;
            14'h1354: rddata <= 8'h7A; 14'h1355: rddata <= 8'h1F; 14'h1356: rddata <= 8'h57; 14'h1357: rddata <= 8'h7B;
            14'h1358: rddata <= 8'h1F; 14'h1359: rddata <= 8'h5F; 14'h135A: rddata <= 8'h78; 14'h135B: rddata <= 8'h1F;
            14'h135C: rddata <= 8'h47; 14'h135D: rddata <= 8'h18; 14'h135E: rddata <= 8'hEF; 14'h135F: rddata <= 8'h00;
            14'h1360: rddata <= 8'h00; 14'h1361: rddata <= 8'h00; 14'h1362: rddata <= 8'h81; 14'h1363: rddata <= 8'h04;
            14'h1364: rddata <= 8'h9A; 14'h1365: rddata <= 8'hF7; 14'h1366: rddata <= 8'h19; 14'h1367: rddata <= 8'h83;
            14'h1368: rddata <= 8'h24; 14'h1369: rddata <= 8'h63; 14'h136A: rddata <= 8'h43; 14'h136B: rddata <= 8'h83;
            14'h136C: rddata <= 8'h75; 14'h136D: rddata <= 8'hCD; 14'h136E: rddata <= 8'h8D; 14'h136F: rddata <= 8'h84;
            14'h1370: rddata <= 8'hA9; 14'h1371: rddata <= 8'h7F; 14'h1372: rddata <= 8'h83; 14'h1373: rddata <= 8'h82;
            14'h1374: rddata <= 8'h04; 14'h1375: rddata <= 8'h00; 14'h1376: rddata <= 8'h00; 14'h1377: rddata <= 8'h00;
            14'h1378: rddata <= 8'h81; 14'h1379: rddata <= 8'hE2; 14'h137A: rddata <= 8'hB0; 14'h137B: rddata <= 8'h4D;
            14'h137C: rddata <= 8'h83; 14'h137D: rddata <= 8'h0A; 14'h137E: rddata <= 8'h72; 14'h137F: rddata <= 8'h11;
            14'h1380: rddata <= 8'h83; 14'h1381: rddata <= 8'hF4; 14'h1382: rddata <= 8'h04; 14'h1383: rddata <= 8'h35;
            14'h1384: rddata <= 8'h7F; 14'h1385: rddata <= 8'hEF; 14'h1386: rddata <= 8'hB7; 14'h1387: rddata <= 8'hEA;
            14'h1388: rddata <= 8'h97; 14'h1389: rddata <= 8'h06; 14'h138A: rddata <= 8'hCD; 14'h138B: rddata <= 8'h95;
            14'h138C: rddata <= 8'h13; 14'h138D: rddata <= 8'h01; 14'h138E: rddata <= 8'h31; 14'h138F: rddata <= 8'h80;
            14'h1390: rddata <= 8'h11; 14'h1391: rddata <= 8'h18; 14'h1392: rddata <= 8'h72; 14'h1393: rddata <= 8'h18;
            14'h1394: rddata <= 8'h36; 14'h1395: rddata <= 8'hCD; 14'h1396: rddata <= 8'h2E; 14'h1397: rddata <= 8'h15;
            14'h1398: rddata <= 8'h3E; 14'h1399: rddata <= 8'h80; 14'h139A: rddata <= 8'h32; 14'h139B: rddata <= 8'hE7;
            14'h139C: rddata <= 8'h38; 14'h139D: rddata <= 8'hA8; 14'h139E: rddata <= 8'hF5; 14'h139F: rddata <= 8'hCD;
            14'h13A0: rddata <= 8'h13; 14'h13A1: rddata <= 8'h15; 14'h13A2: rddata <= 8'h21; 14'h13A3: rddata <= 8'h63;
            14'h13A4: rddata <= 8'h13; 14'h13A5: rddata <= 8'hCD; 14'h13A6: rddata <= 8'h46; 14'h13A7: rddata <= 8'h18;
            14'h13A8: rddata <= 8'hC1; 14'h13A9: rddata <= 8'hE1; 14'h13AA: rddata <= 8'hCD; 14'h13AB: rddata <= 8'h13;
            14'h13AC: rddata <= 8'h15; 14'h13AD: rddata <= 8'hEB; 14'h13AE: rddata <= 8'hCD; 14'h13AF: rddata <= 8'h23;
            14'h13B0: rddata <= 8'h15; 14'h13B1: rddata <= 8'h21; 14'h13B2: rddata <= 8'h74; 14'h13B3: rddata <= 8'h13;
            14'h13B4: rddata <= 8'hCD; 14'h13B5: rddata <= 8'h46; 14'h13B6: rddata <= 8'h18; 14'h13B7: rddata <= 8'hC1;
            14'h13B8: rddata <= 8'hD1; 14'h13B9: rddata <= 8'hCD; 14'h13BA: rddata <= 8'h2F; 14'h13BB: rddata <= 8'h14;
            14'h13BC: rddata <= 8'hF1; 14'h13BD: rddata <= 8'hCD; 14'h13BE: rddata <= 8'h13; 14'h13BF: rddata <= 8'h15;
            14'h13C0: rddata <= 8'hCD; 14'h13C1: rddata <= 8'hF6; 14'h13C2: rddata <= 8'h14; 14'h13C3: rddata <= 8'hC1;
            14'h13C4: rddata <= 8'hD1; 14'h13C5: rddata <= 8'hC3; 14'h13C6: rddata <= 8'h61; 14'h13C7: rddata <= 8'h12;
            14'h13C8: rddata <= 8'h21; 14'h13C9: rddata <= 8'hC1; 14'h13CA: rddata <= 8'hD1; 14'h13CB: rddata <= 8'hEF;
            14'h13CC: rddata <= 8'hC8; 14'h13CD: rddata <= 8'h2E; 14'h13CE: rddata <= 8'h00; 14'h13CF: rddata <= 8'hCD;
            14'h13D0: rddata <= 8'hAC; 14'h13D1: rddata <= 8'h14; 14'h13D2: rddata <= 8'h79; 14'h13D3: rddata <= 8'h32;
            14'h13D4: rddata <= 8'hF6; 14'h13D5: rddata <= 8'h38; 14'h13D6: rddata <= 8'hEB; 14'h13D7: rddata <= 8'h22;
            14'h13D8: rddata <= 8'hF7; 14'h13D9: rddata <= 8'h38; 14'h13DA: rddata <= 8'h01; 14'h13DB: rddata <= 8'h00;
            14'h13DC: rddata <= 8'h00; 14'h13DD: rddata <= 8'h50; 14'h13DE: rddata <= 8'h58; 14'h13DF: rddata <= 8'h21;
            14'h13E0: rddata <= 8'hB0; 14'h13E1: rddata <= 8'h12; 14'h13E2: rddata <= 8'hE5; 14'h13E3: rddata <= 8'h21;
            14'h13E4: rddata <= 8'hEB; 14'h13E5: rddata <= 8'h13; 14'h13E6: rddata <= 8'hE5; 14'h13E7: rddata <= 8'hE5;
            14'h13E8: rddata <= 8'h21; 14'h13E9: rddata <= 8'hE4; 14'h13EA: rddata <= 8'h38; 14'h13EB: rddata <= 8'h7E;
            14'h13EC: rddata <= 8'h23; 14'h13ED: rddata <= 8'hB7; 14'h13EE: rddata <= 8'h28; 14'h13EF: rddata <= 8'h2C;
            14'h13F0: rddata <= 8'hE5; 14'h13F1: rddata <= 8'h2E; 14'h13F2: rddata <= 8'h08; 14'h13F3: rddata <= 8'h1F;
            14'h13F4: rddata <= 8'h67; 14'h13F5: rddata <= 8'h79; 14'h13F6: rddata <= 8'h30; 14'h13F7: rddata <= 8'h0B;
            14'h13F8: rddata <= 8'hE5; 14'h13F9: rddata <= 8'h2A; 14'h13FA: rddata <= 8'hF7; 14'h13FB: rddata <= 8'h38;
            14'h13FC: rddata <= 8'h19; 14'h13FD: rddata <= 8'hEB; 14'h13FE: rddata <= 8'hE1; 14'h13FF: rddata <= 8'h3A;
            14'h1400: rddata <= 8'hF6; 14'h1401: rddata <= 8'h38; 14'h1402: rddata <= 8'h89; 14'h1403: rddata <= 8'h1F;
            14'h1404: rddata <= 8'h4F; 14'h1405: rddata <= 8'h7A; 14'h1406: rddata <= 8'h1F; 14'h1407: rddata <= 8'h57;
            14'h1408: rddata <= 8'h7B; 14'h1409: rddata <= 8'h1F; 14'h140A: rddata <= 8'h5F; 14'h140B: rddata <= 8'h78;
            14'h140C: rddata <= 8'h1F; 14'h140D: rddata <= 8'h47; 14'h140E: rddata <= 8'hE6; 14'h140F: rddata <= 8'h10;
            14'h1410: rddata <= 8'h28; 14'h1411: rddata <= 8'h04; 14'h1412: rddata <= 8'h78; 14'h1413: rddata <= 8'hF6;
            14'h1414: rddata <= 8'h20; 14'h1415: rddata <= 8'h47; 14'h1416: rddata <= 8'h2D; 14'h1417: rddata <= 8'h7C;
            14'h1418: rddata <= 8'h20; 14'h1419: rddata <= 8'hD9; 14'h141A: rddata <= 8'hE1; 14'h141B: rddata <= 8'hC9;
            14'h141C: rddata <= 8'h43; 14'h141D: rddata <= 8'h5A; 14'h141E: rddata <= 8'h51; 14'h141F: rddata <= 8'h4F;
            14'h1420: rddata <= 8'hC9; 14'h1421: rddata <= 8'hCD; 14'h1422: rddata <= 8'h13; 14'h1423: rddata <= 8'h15;
            14'h1424: rddata <= 8'h01; 14'h1425: rddata <= 8'h20; 14'h1426: rddata <= 8'h84; 14'h1427: rddata <= 8'h11;
            14'h1428: rddata <= 8'h00; 14'h1429: rddata <= 8'h00; 14'h142A: rddata <= 8'hCD; 14'h142B: rddata <= 8'h23;
            14'h142C: rddata <= 8'h15; 14'h142D: rddata <= 8'hC1; 14'h142E: rddata <= 8'hD1; 14'h142F: rddata <= 8'hEF;
            14'h1430: rddata <= 8'hCA; 14'h1431: rddata <= 8'hC7; 14'h1432: rddata <= 8'h03; 14'h1433: rddata <= 8'h2E;
            14'h1434: rddata <= 8'hFF; 14'h1435: rddata <= 8'hCD; 14'h1436: rddata <= 8'hAC; 14'h1437: rddata <= 8'h14;
            14'h1438: rddata <= 8'h34; 14'h1439: rddata <= 8'hCA; 14'h143A: rddata <= 8'hD3; 14'h143B: rddata <= 8'h03;
            14'h143C: rddata <= 8'h34; 14'h143D: rddata <= 8'hCA; 14'h143E: rddata <= 8'hD3; 14'h143F: rddata <= 8'h03;
            14'h1440: rddata <= 8'h2B; 14'h1441: rddata <= 8'h7E; 14'h1442: rddata <= 8'h32; 14'h1443: rddata <= 8'h19;
            14'h1444: rddata <= 8'h38; 14'h1445: rddata <= 8'h2B; 14'h1446: rddata <= 8'h7E; 14'h1447: rddata <= 8'h32;
            14'h1448: rddata <= 8'h15; 14'h1449: rddata <= 8'h38; 14'h144A: rddata <= 8'h2B; 14'h144B: rddata <= 8'h7E;
            14'h144C: rddata <= 8'h32; 14'h144D: rddata <= 8'h11; 14'h144E: rddata <= 8'h38; 14'h144F: rddata <= 8'h41;
            14'h1450: rddata <= 8'hEB; 14'h1451: rddata <= 8'hAF; 14'h1452: rddata <= 8'h4F; 14'h1453: rddata <= 8'h57;
            14'h1454: rddata <= 8'h5F; 14'h1455: rddata <= 8'h32; 14'h1456: rddata <= 8'h1C; 14'h1457: rddata <= 8'h38;
            14'h1458: rddata <= 8'hE5; 14'h1459: rddata <= 8'hC5; 14'h145A: rddata <= 8'h7D; 14'h145B: rddata <= 8'hCD;
            14'h145C: rddata <= 8'h10; 14'h145D: rddata <= 8'h38; 14'h145E: rddata <= 8'hDE; 14'h145F: rddata <= 8'h00;
            14'h1460: rddata <= 8'h3F; 14'h1461: rddata <= 8'h30; 14'h1462: rddata <= 8'h07; 14'h1463: rddata <= 8'h32;
            14'h1464: rddata <= 8'h1C; 14'h1465: rddata <= 8'h38; 14'h1466: rddata <= 8'hF1; 14'h1467: rddata <= 8'hF1;
            14'h1468: rddata <= 8'h37; 14'h1469: rddata <= 8'hD2; 14'h146A: rddata <= 8'hC1; 14'h146B: rddata <= 8'hE1;
            14'h146C: rddata <= 8'h79; 14'h146D: rddata <= 8'h3C; 14'h146E: rddata <= 8'h3D; 14'h146F: rddata <= 8'h1F;
            14'h1470: rddata <= 8'hF2; 14'h1471: rddata <= 8'h87; 14'h1472: rddata <= 8'h14; 14'h1473: rddata <= 8'h17;
            14'h1474: rddata <= 8'h3A; 14'h1475: rddata <= 8'h1C; 14'h1476: rddata <= 8'h38; 14'h1477: rddata <= 8'h1F;
            14'h1478: rddata <= 8'hE6; 14'h1479: rddata <= 8'hC0; 14'h147A: rddata <= 8'hF5; 14'h147B: rddata <= 8'h78;
            14'h147C: rddata <= 8'hB4; 14'h147D: rddata <= 8'hB5; 14'h147E: rddata <= 8'h28; 14'h147F: rddata <= 8'h02;
            14'h1480: rddata <= 8'h3E; 14'h1481: rddata <= 8'h20; 14'h1482: rddata <= 8'hE1; 14'h1483: rddata <= 8'hB4;
            14'h1484: rddata <= 8'hC3; 14'h1485: rddata <= 8'hF2; 14'h1486: rddata <= 8'h12; 14'h1487: rddata <= 8'h17;
            14'h1488: rddata <= 8'h7B; 14'h1489: rddata <= 8'h17; 14'h148A: rddata <= 8'h5F; 14'h148B: rddata <= 8'h7A;
            14'h148C: rddata <= 8'h17; 14'h148D: rddata <= 8'h57; 14'h148E: rddata <= 8'h79; 14'h148F: rddata <= 8'h17;
            14'h1490: rddata <= 8'h4F; 14'h1491: rddata <= 8'h29; 14'h1492: rddata <= 8'h78; 14'h1493: rddata <= 8'h17;
            14'h1494: rddata <= 8'h47; 14'h1495: rddata <= 8'h3A; 14'h1496: rddata <= 8'h1C; 14'h1497: rddata <= 8'h38;
            14'h1498: rddata <= 8'h17; 14'h1499: rddata <= 8'h32; 14'h149A: rddata <= 8'h1C; 14'h149B: rddata <= 8'h38;
            14'h149C: rddata <= 8'h79; 14'h149D: rddata <= 8'hB2; 14'h149E: rddata <= 8'hB3; 14'h149F: rddata <= 8'h20;
            14'h14A0: rddata <= 8'hB7; 14'h14A1: rddata <= 8'hE5; 14'h14A2: rddata <= 8'h21; 14'h14A3: rddata <= 8'hE7;
            14'h14A4: rddata <= 8'h38; 14'h14A5: rddata <= 8'h35; 14'h14A6: rddata <= 8'hE1; 14'h14A7: rddata <= 8'h20;
            14'h14A8: rddata <= 8'hAF; 14'h14A9: rddata <= 8'hC3; 14'h14AA: rddata <= 8'hC3; 14'h14AB: rddata <= 8'h12;
            14'h14AC: rddata <= 8'h78; 14'h14AD: rddata <= 8'hB7; 14'h14AE: rddata <= 8'h28; 14'h14AF: rddata <= 8'h1D;
            14'h14B0: rddata <= 8'h7D; 14'h14B1: rddata <= 8'h21; 14'h14B2: rddata <= 8'hE7; 14'h14B3: rddata <= 8'h38;
            14'h14B4: rddata <= 8'hAE; 14'h14B5: rddata <= 8'h80; 14'h14B6: rddata <= 8'h47; 14'h14B7: rddata <= 8'h1F;
            14'h14B8: rddata <= 8'hA8; 14'h14B9: rddata <= 8'h78; 14'h14BA: rddata <= 8'hF2; 14'h14BB: rddata <= 8'hCC;
            14'h14BC: rddata <= 8'h14; 14'h14BD: rddata <= 8'hC6; 14'h14BE: rddata <= 8'h80; 14'h14BF: rddata <= 8'h77;
            14'h14C0: rddata <= 8'hCA; 14'h14C1: rddata <= 8'h1A; 14'h14C2: rddata <= 8'h14; 14'h14C3: rddata <= 8'hCD;
            14'h14C4: rddata <= 8'h46; 14'h14C5: rddata <= 8'h15; 14'h14C6: rddata <= 8'h77; 14'h14C7: rddata <= 8'h2B;
            14'h14C8: rddata <= 8'hC9; 14'h14C9: rddata <= 8'hEF; 14'h14CA: rddata <= 8'h2F; 14'h14CB: rddata <= 8'hE1;
            14'h14CC: rddata <= 8'hB7; 14'h14CD: rddata <= 8'hE1; 14'h14CE: rddata <= 8'hF2; 14'h14CF: rddata <= 8'hC3;
            14'h14D0: rddata <= 8'h12; 14'h14D1: rddata <= 8'hC3; 14'h14D2: rddata <= 8'hD3; 14'h14D3: rddata <= 8'h03;
            14'h14D4: rddata <= 8'hCD; 14'h14D5: rddata <= 8'h2E; 14'h14D6: rddata <= 8'h15; 14'h14D7: rddata <= 8'h78;
            14'h14D8: rddata <= 8'hB7; 14'h14D9: rddata <= 8'hC8; 14'h14DA: rddata <= 8'hC6; 14'h14DB: rddata <= 8'h02;
            14'h14DC: rddata <= 8'hDA; 14'h14DD: rddata <= 8'hD3; 14'h14DE: rddata <= 8'h03; 14'h14DF: rddata <= 8'h47;
            14'h14E0: rddata <= 8'hCD; 14'h14E1: rddata <= 8'h61; 14'h14E2: rddata <= 8'h12; 14'h14E3: rddata <= 8'h21;
            14'h14E4: rddata <= 8'hE7; 14'h14E5: rddata <= 8'h38; 14'h14E6: rddata <= 8'h34; 14'h14E7: rddata <= 8'hC0;
            14'h14E8: rddata <= 8'hC3; 14'h14E9: rddata <= 8'hD3; 14'h14EA: rddata <= 8'h03; 14'h14EB: rddata <= 8'h3A;
            14'h14EC: rddata <= 8'hE6; 14'h14ED: rddata <= 8'h38; 14'h14EE: rddata <= 8'hFE; 14'h14EF: rddata <= 8'h2F;
            14'h14F0: rddata <= 8'h17; 14'h14F1: rddata <= 8'h9F; 14'h14F2: rddata <= 8'hC0; 14'h14F3: rddata <= 8'h3C;
            14'h14F4: rddata <= 8'hC9; 14'h14F5: rddata <= 8'hEF; 14'h14F6: rddata <= 8'h06; 14'h14F7: rddata <= 8'h88;
            14'h14F8: rddata <= 8'h11; 14'h14F9: rddata <= 8'h00; 14'h14FA: rddata <= 8'h00; 14'h14FB: rddata <= 8'h21;
            14'h14FC: rddata <= 8'hE7; 14'h14FD: rddata <= 8'h38; 14'h14FE: rddata <= 8'h4F; 14'h14FF: rddata <= 8'h70;
            14'h1500: rddata <= 8'h06; 14'h1501: rddata <= 8'h00; 14'h1502: rddata <= 8'h23; 14'h1503: rddata <= 8'h36;
            14'h1504: rddata <= 8'h80; 14'h1505: rddata <= 8'h17; 14'h1506: rddata <= 8'hC3; 14'h1507: rddata <= 8'hAD;
            14'h1508: rddata <= 8'h12; 14'h1509: rddata <= 8'hEF; 14'h150A: rddata <= 8'hF0; 14'h150B: rddata <= 8'h21;
            14'h150C: rddata <= 8'hE6; 14'h150D: rddata <= 8'h38; 14'h150E: rddata <= 8'h7E; 14'h150F: rddata <= 8'hEE;
            14'h1510: rddata <= 8'h80; 14'h1511: rddata <= 8'h77; 14'h1512: rddata <= 8'hC9; 14'h1513: rddata <= 8'hEB;
            14'h1514: rddata <= 8'h2A; 14'h1515: rddata <= 8'hE4; 14'h1516: rddata <= 8'h38; 14'h1517: rddata <= 8'hE3;
            14'h1518: rddata <= 8'hE5; 14'h1519: rddata <= 8'h2A; 14'h151A: rddata <= 8'hE6; 14'h151B: rddata <= 8'h38;
            14'h151C: rddata <= 8'hE3; 14'h151D: rddata <= 8'hE5; 14'h151E: rddata <= 8'hEB; 14'h151F: rddata <= 8'hC9;
            14'h1520: rddata <= 8'hCD; 14'h1521: rddata <= 8'h31; 14'h1522: rddata <= 8'h15; 14'h1523: rddata <= 8'hEB;
            14'h1524: rddata <= 8'h22; 14'h1525: rddata <= 8'hE4; 14'h1526: rddata <= 8'h38; 14'h1527: rddata <= 8'h60;
            14'h1528: rddata <= 8'h69; 14'h1529: rddata <= 8'h22; 14'h152A: rddata <= 8'hE6; 14'h152B: rddata <= 8'h38;
            14'h152C: rddata <= 8'hEB; 14'h152D: rddata <= 8'hC9; 14'h152E: rddata <= 8'h21; 14'h152F: rddata <= 8'hE4;
            14'h1530: rddata <= 8'h38; 14'h1531: rddata <= 8'h5E; 14'h1532: rddata <= 8'h23; 14'h1533: rddata <= 8'h56;
            14'h1534: rddata <= 8'h23; 14'h1535: rddata <= 8'h4E; 14'h1536: rddata <= 8'h23; 14'h1537: rddata <= 8'h46;
            14'h1538: rddata <= 8'h23; 14'h1539: rddata <= 8'hC9; 14'h153A: rddata <= 8'h11; 14'h153B: rddata <= 8'hE4;
            14'h153C: rddata <= 8'h38; 14'h153D: rddata <= 8'h06; 14'h153E: rddata <= 8'h04; 14'h153F: rddata <= 8'h1A;
            14'h1540: rddata <= 8'h77; 14'h1541: rddata <= 8'h13; 14'h1542: rddata <= 8'h23; 14'h1543: rddata <= 8'h10;
            14'h1544: rddata <= 8'hFA; 14'h1545: rddata <= 8'hC9; 14'h1546: rddata <= 8'h21; 14'h1547: rddata <= 8'hE6;
            14'h1548: rddata <= 8'h38; 14'h1549: rddata <= 8'h7E; 14'h154A: rddata <= 8'h07; 14'h154B: rddata <= 8'h37;
            14'h154C: rddata <= 8'h1F; 14'h154D: rddata <= 8'h77; 14'h154E: rddata <= 8'h3F; 14'h154F: rddata <= 8'h1F;
            14'h1550: rddata <= 8'h23; 14'h1551: rddata <= 8'h23; 14'h1552: rddata <= 8'h77; 14'h1553: rddata <= 8'h79;
            14'h1554: rddata <= 8'h07; 14'h1555: rddata <= 8'h37; 14'h1556: rddata <= 8'h1F; 14'h1557: rddata <= 8'h4F;
            14'h1558: rddata <= 8'h1F; 14'h1559: rddata <= 8'hAE; 14'h155A: rddata <= 8'hC9; 14'h155B: rddata <= 8'h78;
            14'h155C: rddata <= 8'hB7; 14'h155D: rddata <= 8'hCA; 14'h155E: rddata <= 8'h28; 14'h155F: rddata <= 8'h00;
            14'h1560: rddata <= 8'h21; 14'h1561: rddata <= 8'hEF; 14'h1562: rddata <= 8'h14; 14'h1563: rddata <= 8'hE5;
            14'h1564: rddata <= 8'hEF; 14'h1565: rddata <= 8'h79; 14'h1566: rddata <= 8'hC8; 14'h1567: rddata <= 8'h21;
            14'h1568: rddata <= 8'hE6; 14'h1569: rddata <= 8'h38; 14'h156A: rddata <= 8'hAE; 14'h156B: rddata <= 8'h79;
            14'h156C: rddata <= 8'hF8; 14'h156D: rddata <= 8'hCD; 14'h156E: rddata <= 8'h73; 14'h156F: rddata <= 8'h15;
            14'h1570: rddata <= 8'h1F; 14'h1571: rddata <= 8'hA9; 14'h1572: rddata <= 8'hC9; 14'h1573: rddata <= 8'h23;
            14'h1574: rddata <= 8'h78; 14'h1575: rddata <= 8'hBE; 14'h1576: rddata <= 8'hC0; 14'h1577: rddata <= 8'h2B;
            14'h1578: rddata <= 8'h79; 14'h1579: rddata <= 8'hBE; 14'h157A: rddata <= 8'hC0; 14'h157B: rddata <= 8'h2B;
            14'h157C: rddata <= 8'h7A; 14'h157D: rddata <= 8'hBE; 14'h157E: rddata <= 8'hC0; 14'h157F: rddata <= 8'h2B;
            14'h1580: rddata <= 8'h7B; 14'h1581: rddata <= 8'h96; 14'h1582: rddata <= 8'hC0; 14'h1583: rddata <= 8'hE1;
            14'h1584: rddata <= 8'hE1; 14'h1585: rddata <= 8'hC9; 14'h1586: rddata <= 8'h47; 14'h1587: rddata <= 8'h4F;
            14'h1588: rddata <= 8'h57; 14'h1589: rddata <= 8'h5F; 14'h158A: rddata <= 8'hB7; 14'h158B: rddata <= 8'hC8;
            14'h158C: rddata <= 8'hE5; 14'h158D: rddata <= 8'hCD; 14'h158E: rddata <= 8'h2E; 14'h158F: rddata <= 8'h15;
            14'h1590: rddata <= 8'hCD; 14'h1591: rddata <= 8'h46; 14'h1592: rddata <= 8'h15; 14'h1593: rddata <= 8'hAE;
            14'h1594: rddata <= 8'h67; 14'h1595: rddata <= 8'hFC; 14'h1596: rddata <= 8'hAA; 14'h1597: rddata <= 8'h15;
            14'h1598: rddata <= 8'h3E; 14'h1599: rddata <= 8'h98; 14'h159A: rddata <= 8'h90; 14'h159B: rddata <= 8'hCD;
            14'h159C: rddata <= 8'h30; 14'h159D: rddata <= 8'h13; 14'h159E: rddata <= 8'h7C; 14'h159F: rddata <= 8'h17;
            14'h15A0: rddata <= 8'hDC; 14'h15A1: rddata <= 8'h03; 14'h15A2: rddata <= 8'h13; 14'h15A3: rddata <= 8'h06;
            14'h15A4: rddata <= 8'h00; 14'h15A5: rddata <= 8'hDC; 14'h15A6: rddata <= 8'h1C; 14'h15A7: rddata <= 8'h13;
            14'h15A8: rddata <= 8'hE1; 14'h15A9: rddata <= 8'hC9; 14'h15AA: rddata <= 8'h1B; 14'h15AB: rddata <= 8'h7A;
            14'h15AC: rddata <= 8'hA3; 14'h15AD: rddata <= 8'h3C; 14'h15AE: rddata <= 8'hC0; 14'h15AF: rddata <= 8'h0B;
            14'h15B0: rddata <= 8'hC9; 14'h15B1: rddata <= 8'h21; 14'h15B2: rddata <= 8'hE7; 14'h15B3: rddata <= 8'h38;
            14'h15B4: rddata <= 8'h7E; 14'h15B5: rddata <= 8'hFE; 14'h15B6: rddata <= 8'h98; 14'h15B7: rddata <= 8'h3A;
            14'h15B8: rddata <= 8'hE4; 14'h15B9: rddata <= 8'h38; 14'h15BA: rddata <= 8'hD0; 14'h15BB: rddata <= 8'h7E;
            14'h15BC: rddata <= 8'hCD; 14'h15BD: rddata <= 8'h86; 14'h15BE: rddata <= 8'h15; 14'h15BF: rddata <= 8'h36;
            14'h15C0: rddata <= 8'h98; 14'h15C1: rddata <= 8'h7B; 14'h15C2: rddata <= 8'hF5; 14'h15C3: rddata <= 8'h79;
            14'h15C4: rddata <= 8'h17; 14'h15C5: rddata <= 8'hCD; 14'h15C6: rddata <= 8'hAD; 14'h15C7: rddata <= 8'h12;
            14'h15C8: rddata <= 8'hF1; 14'h15C9: rddata <= 8'hC9; 14'h15CA: rddata <= 8'h21; 14'h15CB: rddata <= 8'h00;
            14'h15CC: rddata <= 8'h00; 14'h15CD: rddata <= 8'h78; 14'h15CE: rddata <= 8'hB1; 14'h15CF: rddata <= 8'hC8;
            14'h15D0: rddata <= 8'h3E; 14'h15D1: rddata <= 8'h10; 14'h15D2: rddata <= 8'h29; 14'h15D3: rddata <= 8'hDA;
            14'h15D4: rddata <= 8'hCD; 14'h15D5: rddata <= 8'h11; 14'h15D6: rddata <= 8'hEB; 14'h15D7: rddata <= 8'h29;
            14'h15D8: rddata <= 8'hEB; 14'h15D9: rddata <= 8'hD2; 14'h15DA: rddata <= 8'hE0; 14'h15DB: rddata <= 8'h15;
            14'h15DC: rddata <= 8'h09; 14'h15DD: rddata <= 8'hDA; 14'h15DE: rddata <= 8'hCD; 14'h15DF: rddata <= 8'h11;
            14'h15E0: rddata <= 8'h3D; 14'h15E1: rddata <= 8'hC2; 14'h15E2: rddata <= 8'hD2; 14'h15E3: rddata <= 8'h15;
            14'h15E4: rddata <= 8'hC9; 14'h15E5: rddata <= 8'hFE; 14'h15E6: rddata <= 8'h2D; 14'h15E7: rddata <= 8'hF5;
            14'h15E8: rddata <= 8'h28; 14'h15E9: rddata <= 8'h05; 14'h15EA: rddata <= 8'hFE; 14'h15EB: rddata <= 8'h2B;
            14'h15EC: rddata <= 8'h28; 14'h15ED: rddata <= 8'h01; 14'h15EE: rddata <= 8'h2B; 14'h15EF: rddata <= 8'hCD;
            14'h15F0: rddata <= 8'hC3; 14'h15F1: rddata <= 8'h12; 14'h15F2: rddata <= 8'h47; 14'h15F3: rddata <= 8'h57;
            14'h15F4: rddata <= 8'h5F; 14'h15F5: rddata <= 8'h2F; 14'h15F6: rddata <= 8'h4F; 14'h15F7: rddata <= 8'hD7;
            14'h15F8: rddata <= 8'hDA; 14'h15F9: rddata <= 8'h3F; 14'h15FA: rddata <= 8'h16; 14'h15FB: rddata <= 8'hFE;
            14'h15FC: rddata <= 8'h2E; 14'h15FD: rddata <= 8'hCA; 14'h15FE: rddata <= 8'h1A; 14'h15FF: rddata <= 8'h16;
            14'h1600: rddata <= 8'hFE; 14'h1601: rddata <= 8'h65; 14'h1602: rddata <= 8'hCA; 14'h1603: rddata <= 8'h0A;
            14'h1604: rddata <= 8'h16; 14'h1605: rddata <= 8'hFE; 14'h1606: rddata <= 8'h45; 14'h1607: rddata <= 8'hC2;
            14'h1608: rddata <= 8'h1E; 14'h1609: rddata <= 8'h16; 14'h160A: rddata <= 8'hD7; 14'h160B: rddata <= 8'hCD;
            14'h160C: rddata <= 8'h98; 14'h160D: rddata <= 8'h0A; 14'h160E: rddata <= 8'hD7; 14'h160F: rddata <= 8'hDA;
            14'h1610: rddata <= 8'h61; 14'h1611: rddata <= 8'h16; 14'h1612: rddata <= 8'h14; 14'h1613: rddata <= 8'hC2;
            14'h1614: rddata <= 8'h1E; 14'h1615: rddata <= 8'h16; 14'h1616: rddata <= 8'hAF; 14'h1617: rddata <= 8'h93;
            14'h1618: rddata <= 8'h5F; 14'h1619: rddata <= 8'h0C; 14'h161A: rddata <= 8'h0C; 14'h161B: rddata <= 8'hCA;
            14'h161C: rddata <= 8'hF7; 14'h161D: rddata <= 8'h15; 14'h161E: rddata <= 8'hE5; 14'h161F: rddata <= 8'h7B;
            14'h1620: rddata <= 8'h90; 14'h1621: rddata <= 8'hF4; 14'h1622: rddata <= 8'h37; 14'h1623: rddata <= 8'h16;
            14'h1624: rddata <= 8'hF2; 14'h1625: rddata <= 8'h2D; 14'h1626: rddata <= 8'h16; 14'h1627: rddata <= 8'hF5;
            14'h1628: rddata <= 8'hCD; 14'h1629: rddata <= 8'h21; 14'h162A: rddata <= 8'h14; 14'h162B: rddata <= 8'hF1;
            14'h162C: rddata <= 8'h3C; 14'h162D: rddata <= 8'hC2; 14'h162E: rddata <= 8'h21; 14'h162F: rddata <= 8'h16;
            14'h1630: rddata <= 8'hD1; 14'h1631: rddata <= 8'hF1; 14'h1632: rddata <= 8'hCC; 14'h1633: rddata <= 8'h0B;
            14'h1634: rddata <= 8'h15; 14'h1635: rddata <= 8'hEB; 14'h1636: rddata <= 8'hC9; 14'h1637: rddata <= 8'hC8;
            14'h1638: rddata <= 8'hF5; 14'h1639: rddata <= 8'hCD; 14'h163A: rddata <= 8'hD4; 14'h163B: rddata <= 8'h14;
            14'h163C: rddata <= 8'hF1; 14'h163D: rddata <= 8'h3D; 14'h163E: rddata <= 8'hC9; 14'h163F: rddata <= 8'hD5;
            14'h1640: rddata <= 8'h57; 14'h1641: rddata <= 8'h78; 14'h1642: rddata <= 8'h89; 14'h1643: rddata <= 8'h47;
            14'h1644: rddata <= 8'hC5; 14'h1645: rddata <= 8'hE5; 14'h1646: rddata <= 8'hD5; 14'h1647: rddata <= 8'hCD;
            14'h1648: rddata <= 8'hD4; 14'h1649: rddata <= 8'h14; 14'h164A: rddata <= 8'hF1; 14'h164B: rddata <= 8'hD6;
            14'h164C: rddata <= 8'h30; 14'h164D: rddata <= 8'hCD; 14'h164E: rddata <= 8'h56; 14'h164F: rddata <= 8'h16;
            14'h1650: rddata <= 8'hE1; 14'h1651: rddata <= 8'hC1; 14'h1652: rddata <= 8'hD1; 14'h1653: rddata <= 8'hC3;
            14'h1654: rddata <= 8'hF7; 14'h1655: rddata <= 8'h15; 14'h1656: rddata <= 8'hCD; 14'h1657: rddata <= 8'h13;
            14'h1658: rddata <= 8'h15; 14'h1659: rddata <= 8'hCD; 14'h165A: rddata <= 8'hF6; 14'h165B: rddata <= 8'h14;
            14'h165C: rddata <= 8'hC1; 14'h165D: rddata <= 8'hD1; 14'h165E: rddata <= 8'hC3; 14'h165F: rddata <= 8'h61;
            14'h1660: rddata <= 8'h12; 14'h1661: rddata <= 8'h7B; 14'h1662: rddata <= 8'h07; 14'h1663: rddata <= 8'h07;
            14'h1664: rddata <= 8'h83; 14'h1665: rddata <= 8'h07; 14'h1666: rddata <= 8'h86; 14'h1667: rddata <= 8'hD6;
            14'h1668: rddata <= 8'h30; 14'h1669: rddata <= 8'h5F; 14'h166A: rddata <= 8'hC3; 14'h166B: rddata <= 8'h0E;
            14'h166C: rddata <= 8'h16; 14'h166D: rddata <= 8'hE5; 14'h166E: rddata <= 8'h21; 14'h166F: rddata <= 8'h69;
            14'h1670: rddata <= 8'h03; 14'h1671: rddata <= 8'hCD; 14'h1672: rddata <= 8'h9D; 14'h1673: rddata <= 8'h0E;
            14'h1674: rddata <= 8'hE1; 14'h1675: rddata <= 8'h11; 14'h1676: rddata <= 8'h9C; 14'h1677: rddata <= 8'h0E;
            14'h1678: rddata <= 8'hD5; 14'h1679: rddata <= 8'hEB; 14'h167A: rddata <= 8'hAF; 14'h167B: rddata <= 8'h06;
            14'h167C: rddata <= 8'h98; 14'h167D: rddata <= 8'hCD; 14'h167E: rddata <= 8'hFB; 14'h167F: rddata <= 8'h14;
            14'h1680: rddata <= 8'h21; 14'h1681: rddata <= 8'hE9; 14'h1682: rddata <= 8'h38; 14'h1683: rddata <= 8'hE5;
            14'h1684: rddata <= 8'hEF; 14'h1685: rddata <= 8'h36; 14'h1686: rddata <= 8'h20; 14'h1687: rddata <= 8'hF2;
            14'h1688: rddata <= 8'h8C; 14'h1689: rddata <= 8'h16; 14'h168A: rddata <= 8'h36; 14'h168B: rddata <= 8'h2D;
            14'h168C: rddata <= 8'h23; 14'h168D: rddata <= 8'h36; 14'h168E: rddata <= 8'h30; 14'h168F: rddata <= 8'hCA;
            14'h1690: rddata <= 8'h42; 14'h1691: rddata <= 8'h17; 14'h1692: rddata <= 8'hE5; 14'h1693: rddata <= 8'hFC;
            14'h1694: rddata <= 8'h0B; 14'h1695: rddata <= 8'h15; 14'h1696: rddata <= 8'hAF; 14'h1697: rddata <= 8'hF5;
            14'h1698: rddata <= 8'hCD; 14'h1699: rddata <= 8'h48; 14'h169A: rddata <= 8'h17; 14'h169B: rddata <= 8'h01;
            14'h169C: rddata <= 8'h43; 14'h169D: rddata <= 8'h91; 14'h169E: rddata <= 8'h11; 14'h169F: rddata <= 8'hF8;
            14'h16A0: rddata <= 8'h4F; 14'h16A1: rddata <= 8'hCD; 14'h16A2: rddata <= 8'h5B; 14'h16A3: rddata <= 8'h15;
            14'h16A4: rddata <= 8'hB7; 14'h16A5: rddata <= 8'hE2; 14'h16A6: rddata <= 8'hB9; 14'h16A7: rddata <= 8'h16;
            14'h16A8: rddata <= 8'hF1; 14'h16A9: rddata <= 8'hCD; 14'h16AA: rddata <= 8'h38; 14'h16AB: rddata <= 8'h16;
            14'h16AC: rddata <= 8'hF5; 14'h16AD: rddata <= 8'hC3; 14'h16AE: rddata <= 8'h9B; 14'h16AF: rddata <= 8'h16;
            14'h16B0: rddata <= 8'hCD; 14'h16B1: rddata <= 8'h21; 14'h16B2: rddata <= 8'h14; 14'h16B3: rddata <= 8'hF1;
            14'h16B4: rddata <= 8'h3C; 14'h16B5: rddata <= 8'hF5; 14'h16B6: rddata <= 8'hCD; 14'h16B7: rddata <= 8'h48;
            14'h16B8: rddata <= 8'h17; 14'h16B9: rddata <= 8'hCD; 14'h16BA: rddata <= 8'h50; 14'h16BB: rddata <= 8'h12;
            14'h16BC: rddata <= 8'h3C; 14'h16BD: rddata <= 8'hCD; 14'h16BE: rddata <= 8'h86; 14'h16BF: rddata <= 8'h15;
            14'h16C0: rddata <= 8'hCD; 14'h16C1: rddata <= 8'h23; 14'h16C2: rddata <= 8'h15; 14'h16C3: rddata <= 8'h01;
            14'h16C4: rddata <= 8'h06; 14'h16C5: rddata <= 8'h03; 14'h16C6: rddata <= 8'hF1; 14'h16C7: rddata <= 8'h81;
            14'h16C8: rddata <= 8'h3C; 14'h16C9: rddata <= 8'hFA; 14'h16CA: rddata <= 8'hD5; 14'h16CB: rddata <= 8'h16;
            14'h16CC: rddata <= 8'hFE; 14'h16CD: rddata <= 8'h08; 14'h16CE: rddata <= 8'hD2; 14'h16CF: rddata <= 8'hD5;
            14'h16D0: rddata <= 8'h16; 14'h16D1: rddata <= 8'h3C; 14'h16D2: rddata <= 8'h47; 14'h16D3: rddata <= 8'h3E;
            14'h16D4: rddata <= 8'h02; 14'h16D5: rddata <= 8'h3D; 14'h16D6: rddata <= 8'h3D; 14'h16D7: rddata <= 8'hE1;
            14'h16D8: rddata <= 8'hF5; 14'h16D9: rddata <= 8'h11; 14'h16DA: rddata <= 8'h5E; 14'h16DB: rddata <= 8'h17;
            14'h16DC: rddata <= 8'h05; 14'h16DD: rddata <= 8'hC2; 14'h16DE: rddata <= 8'hE6; 14'h16DF: rddata <= 8'h16;
            14'h16E0: rddata <= 8'h36; 14'h16E1: rddata <= 8'h2E; 14'h16E2: rddata <= 8'h23; 14'h16E3: rddata <= 8'h36;
            14'h16E4: rddata <= 8'h30; 14'h16E5: rddata <= 8'h23; 14'h16E6: rddata <= 8'h05; 14'h16E7: rddata <= 8'h36;
            14'h16E8: rddata <= 8'h2E; 14'h16E9: rddata <= 8'hCC; 14'h16EA: rddata <= 8'h38; 14'h16EB: rddata <= 8'h15;
            14'h16EC: rddata <= 8'hC5; 14'h16ED: rddata <= 8'hE5; 14'h16EE: rddata <= 8'hD5; 14'h16EF: rddata <= 8'hCD;
            14'h16F0: rddata <= 8'h2E; 14'h16F1: rddata <= 8'h15; 14'h16F2: rddata <= 8'hE1; 14'h16F3: rddata <= 8'h06;
            14'h16F4: rddata <= 8'h2F; 14'h16F5: rddata <= 8'h04; 14'h16F6: rddata <= 8'h7B; 14'h16F7: rddata <= 8'h96;
            14'h16F8: rddata <= 8'h5F; 14'h16F9: rddata <= 8'h23; 14'h16FA: rddata <= 8'h7A; 14'h16FB: rddata <= 8'h9E;
            14'h16FC: rddata <= 8'h57; 14'h16FD: rddata <= 8'h23; 14'h16FE: rddata <= 8'h79; 14'h16FF: rddata <= 8'h9E;
            14'h1700: rddata <= 8'h4F; 14'h1701: rddata <= 8'h2B; 14'h1702: rddata <= 8'h2B; 14'h1703: rddata <= 8'hD2;
            14'h1704: rddata <= 8'hF5; 14'h1705: rddata <= 8'h16; 14'h1706: rddata <= 8'hCD; 14'h1707: rddata <= 8'h10;
            14'h1708: rddata <= 8'h13; 14'h1709: rddata <= 8'h23; 14'h170A: rddata <= 8'hCD; 14'h170B: rddata <= 8'h23;
            14'h170C: rddata <= 8'h15; 14'h170D: rddata <= 8'hEB; 14'h170E: rddata <= 8'hE1; 14'h170F: rddata <= 8'h70;
            14'h1710: rddata <= 8'h23; 14'h1711: rddata <= 8'hC1; 14'h1712: rddata <= 8'h0D; 14'h1713: rddata <= 8'hC2;
            14'h1714: rddata <= 8'hE6; 14'h1715: rddata <= 8'h16; 14'h1716: rddata <= 8'h05; 14'h1717: rddata <= 8'hCA;
            14'h1718: rddata <= 8'h26; 14'h1719: rddata <= 8'h17; 14'h171A: rddata <= 8'h2B; 14'h171B: rddata <= 8'h7E;
            14'h171C: rddata <= 8'hFE; 14'h171D: rddata <= 8'h30; 14'h171E: rddata <= 8'hCA; 14'h171F: rddata <= 8'h1A;
            14'h1720: rddata <= 8'h17; 14'h1721: rddata <= 8'hFE; 14'h1722: rddata <= 8'h2E; 14'h1723: rddata <= 8'hC4;
            14'h1724: rddata <= 8'h38; 14'h1725: rddata <= 8'h15; 14'h1726: rddata <= 8'hF1; 14'h1727: rddata <= 8'hCA;
            14'h1728: rddata <= 8'h45; 14'h1729: rddata <= 8'h17; 14'h172A: rddata <= 8'h36; 14'h172B: rddata <= 8'h45;
            14'h172C: rddata <= 8'h23; 14'h172D: rddata <= 8'h36; 14'h172E: rddata <= 8'h2B; 14'h172F: rddata <= 8'hF2;
            14'h1730: rddata <= 8'h36; 14'h1731: rddata <= 8'h17; 14'h1732: rddata <= 8'h36; 14'h1733: rddata <= 8'h2D;
            14'h1734: rddata <= 8'h2F; 14'h1735: rddata <= 8'h3C; 14'h1736: rddata <= 8'h06; 14'h1737: rddata <= 8'h2F;
            14'h1738: rddata <= 8'h04; 14'h1739: rddata <= 8'hD6; 14'h173A: rddata <= 8'h0A; 14'h173B: rddata <= 8'hD2;
            14'h173C: rddata <= 8'h38; 14'h173D: rddata <= 8'h17; 14'h173E: rddata <= 8'hC6; 14'h173F: rddata <= 8'h3A;
            14'h1740: rddata <= 8'h23; 14'h1741: rddata <= 8'h70; 14'h1742: rddata <= 8'h23; 14'h1743: rddata <= 8'h77;
            14'h1744: rddata <= 8'h23; 14'h1745: rddata <= 8'h71; 14'h1746: rddata <= 8'hE1; 14'h1747: rddata <= 8'hC9;
            14'h1748: rddata <= 8'h01; 14'h1749: rddata <= 8'h74; 14'h174A: rddata <= 8'h94; 14'h174B: rddata <= 8'h11;
            14'h174C: rddata <= 8'hF7; 14'h174D: rddata <= 8'h23; 14'h174E: rddata <= 8'hCD; 14'h174F: rddata <= 8'h5B;
            14'h1750: rddata <= 8'h15; 14'h1751: rddata <= 8'hB7; 14'h1752: rddata <= 8'hE1; 14'h1753: rddata <= 8'hE2;
            14'h1754: rddata <= 8'hB0; 14'h1755: rddata <= 8'h16; 14'h1756: rddata <= 8'hE9; 14'h1757: rddata <= 8'h00;
            14'h1758: rddata <= 8'h00; 14'h1759: rddata <= 8'h00; 14'h175A: rddata <= 8'h80; 14'h175B: rddata <= 8'h40;
            14'h175C: rddata <= 8'h42; 14'h175D: rddata <= 8'h0F; 14'h175E: rddata <= 8'hA0; 14'h175F: rddata <= 8'h86;
            14'h1760: rddata <= 8'h01; 14'h1761: rddata <= 8'h10; 14'h1762: rddata <= 8'h27; 14'h1763: rddata <= 8'h00;
            14'h1764: rddata <= 8'hE8; 14'h1765: rddata <= 8'h03; 14'h1766: rddata <= 8'h00; 14'h1767: rddata <= 8'h64;
            14'h1768: rddata <= 8'h00; 14'h1769: rddata <= 8'h00; 14'h176A: rddata <= 8'h0A; 14'h176B: rddata <= 8'h00;
            14'h176C: rddata <= 8'h00; 14'h176D: rddata <= 8'h01; 14'h176E: rddata <= 8'h00; 14'h176F: rddata <= 8'h00;
            14'h1770: rddata <= 8'h21; 14'h1771: rddata <= 8'h0B; 14'h1772: rddata <= 8'h15; 14'h1773: rddata <= 8'hE3;
            14'h1774: rddata <= 8'hE9; 14'h1775: rddata <= 8'hCD; 14'h1776: rddata <= 8'h13; 14'h1777: rddata <= 8'h15;
            14'h1778: rddata <= 8'h21; 14'h1779: rddata <= 8'h57; 14'h177A: rddata <= 8'h17; 14'h177B: rddata <= 8'hCD;
            14'h177C: rddata <= 8'h20; 14'h177D: rddata <= 8'h15; 14'h177E: rddata <= 8'hC1; 14'h177F: rddata <= 8'hD1;
            14'h1780: rddata <= 8'hEF; 14'h1781: rddata <= 8'h78; 14'h1782: rddata <= 8'hCA; 14'h1783: rddata <= 8'hCD;
            14'h1784: rddata <= 8'h17; 14'h1785: rddata <= 8'hF2; 14'h1786: rddata <= 8'h8C; 14'h1787: rddata <= 8'h17;
            14'h1788: rddata <= 8'hB7; 14'h1789: rddata <= 8'hCA; 14'h178A: rddata <= 8'hC7; 14'h178B: rddata <= 8'h03;
            14'h178C: rddata <= 8'hB7; 14'h178D: rddata <= 8'hCA; 14'h178E: rddata <= 8'hC4; 14'h178F: rddata <= 8'h12;
            14'h1790: rddata <= 8'hD5; 14'h1791: rddata <= 8'hC5; 14'h1792: rddata <= 8'h79; 14'h1793: rddata <= 8'hF6;
            14'h1794: rddata <= 8'h7F; 14'h1795: rddata <= 8'hCD; 14'h1796: rddata <= 8'h2E; 14'h1797: rddata <= 8'h15;
            14'h1798: rddata <= 8'hF2; 14'h1799: rddata <= 8'hB5; 14'h179A: rddata <= 8'h17; 14'h179B: rddata <= 8'hF5;
            14'h179C: rddata <= 8'h3A; 14'h179D: rddata <= 8'hE7; 14'h179E: rddata <= 8'h38; 14'h179F: rddata <= 8'hFE;
            14'h17A0: rddata <= 8'h99; 14'h17A1: rddata <= 8'h38; 14'h17A2: rddata <= 8'h03; 14'h17A3: rddata <= 8'hF1;
            14'h17A4: rddata <= 8'h18; 14'h17A5: rddata <= 8'h0F; 14'h17A6: rddata <= 8'hF1; 14'h17A7: rddata <= 8'hD5;
            14'h17A8: rddata <= 8'hC5; 14'h17A9: rddata <= 8'hCD; 14'h17AA: rddata <= 8'hB1; 14'h17AB: rddata <= 8'h15;
            14'h17AC: rddata <= 8'hC1; 14'h17AD: rddata <= 8'hD1; 14'h17AE: rddata <= 8'hF5; 14'h17AF: rddata <= 8'hCD;
            14'h17B0: rddata <= 8'h5B; 14'h17B1: rddata <= 8'h15; 14'h17B2: rddata <= 8'hE1; 14'h17B3: rddata <= 8'h7C;
            14'h17B4: rddata <= 8'h1F; 14'h17B5: rddata <= 8'hE1; 14'h17B6: rddata <= 8'h22; 14'h17B7: rddata <= 8'hE6;
            14'h17B8: rddata <= 8'h38; 14'h17B9: rddata <= 8'hE1; 14'h17BA: rddata <= 8'h22; 14'h17BB: rddata <= 8'hE4;
            14'h17BC: rddata <= 8'h38; 14'h17BD: rddata <= 8'hDC; 14'h17BE: rddata <= 8'h70; 14'h17BF: rddata <= 8'h17;
            14'h17C0: rddata <= 8'hCC; 14'h17C1: rddata <= 8'h0B; 14'h17C2: rddata <= 8'h15; 14'h17C3: rddata <= 8'hD5;
            14'h17C4: rddata <= 8'hC5; 14'h17C5: rddata <= 8'hCD; 14'h17C6: rddata <= 8'h85; 14'h17C7: rddata <= 8'h13;
            14'h17C8: rddata <= 8'hC1; 14'h17C9: rddata <= 8'hD1; 14'h17CA: rddata <= 8'hCD; 14'h17CB: rddata <= 8'hCB;
            14'h17CC: rddata <= 8'h13; 14'h17CD: rddata <= 8'h01; 14'h17CE: rddata <= 8'h38; 14'h17CF: rddata <= 8'h81;
            14'h17D0: rddata <= 8'h11; 14'h17D1: rddata <= 8'h3B; 14'h17D2: rddata <= 8'hAA; 14'h17D3: rddata <= 8'hCD;
            14'h17D4: rddata <= 8'hCB; 14'h17D5: rddata <= 8'h13; 14'h17D6: rddata <= 8'h3A; 14'h17D7: rddata <= 8'hE7;
            14'h17D8: rddata <= 8'h38; 14'h17D9: rddata <= 8'hFE; 14'h17DA: rddata <= 8'h88; 14'h17DB: rddata <= 8'h30;
            14'h17DC: rddata <= 8'h22; 14'h17DD: rddata <= 8'hFE; 14'h17DE: rddata <= 8'h68; 14'h17DF: rddata <= 8'h38;
            14'h17E0: rddata <= 8'h30; 14'h17E1: rddata <= 8'hCD; 14'h17E2: rddata <= 8'h13; 14'h17E3: rddata <= 8'h15;
            14'h17E4: rddata <= 8'hCD; 14'h17E5: rddata <= 8'hB1; 14'h17E6: rddata <= 8'h15; 14'h17E7: rddata <= 8'hC6;
            14'h17E8: rddata <= 8'h81; 14'h17E9: rddata <= 8'hC1; 14'h17EA: rddata <= 8'hD1; 14'h17EB: rddata <= 8'h28;
            14'h17EC: rddata <= 8'h15; 14'h17ED: rddata <= 8'hF5; 14'h17EE: rddata <= 8'hCD; 14'h17EF: rddata <= 8'h5E;
            14'h17F0: rddata <= 8'h12; 14'h17F1: rddata <= 8'h21; 14'h17F2: rddata <= 8'h1A; 14'h17F3: rddata <= 8'h18;
            14'h17F4: rddata <= 8'hCD; 14'h17F5: rddata <= 8'h46; 14'h17F6: rddata <= 8'h18; 14'h17F7: rddata <= 8'hC1;
            14'h17F8: rddata <= 8'h11; 14'h17F9: rddata <= 8'h00; 14'h17FA: rddata <= 8'h00; 14'h17FB: rddata <= 8'h4A;
            14'h17FC: rddata <= 8'hC3; 14'h17FD: rddata <= 8'hCB; 14'h17FE: rddata <= 8'h13; 14'h17FF: rddata <= 8'hCD;
            14'h1800: rddata <= 8'h13; 14'h1801: rddata <= 8'h15; 14'h1802: rddata <= 8'h3A; 14'h1803: rddata <= 8'hE6;
            14'h1804: rddata <= 8'h38; 14'h1805: rddata <= 8'hB7; 14'h1806: rddata <= 8'hF2; 14'h1807: rddata <= 8'h0E;
            14'h1808: rddata <= 8'h18; 14'h1809: rddata <= 8'hF1; 14'h180A: rddata <= 8'hF1; 14'h180B: rddata <= 8'hC3;
            14'h180C: rddata <= 8'hC3; 14'h180D: rddata <= 8'h12; 14'h180E: rddata <= 8'hC3; 14'h180F: rddata <= 8'hD3;
            14'h1810: rddata <= 8'h03; 14'h1811: rddata <= 8'h01; 14'h1812: rddata <= 8'h00; 14'h1813: rddata <= 8'h81;
            14'h1814: rddata <= 8'h11; 14'h1815: rddata <= 8'h00; 14'h1816: rddata <= 8'h00; 14'h1817: rddata <= 8'hC3;
            14'h1818: rddata <= 8'h23; 14'h1819: rddata <= 8'h15; 14'h181A: rddata <= 8'h07; 14'h181B: rddata <= 8'h7C;
            14'h181C: rddata <= 8'h88; 14'h181D: rddata <= 8'h59; 14'h181E: rddata <= 8'h74; 14'h181F: rddata <= 8'hE0;
            14'h1820: rddata <= 8'h97; 14'h1821: rddata <= 8'h26; 14'h1822: rddata <= 8'h77; 14'h1823: rddata <= 8'hC4;
            14'h1824: rddata <= 8'h1D; 14'h1825: rddata <= 8'h1E; 14'h1826: rddata <= 8'h7A; 14'h1827: rddata <= 8'h5E;
            14'h1828: rddata <= 8'h50; 14'h1829: rddata <= 8'h63; 14'h182A: rddata <= 8'h7C; 14'h182B: rddata <= 8'h1A;
            14'h182C: rddata <= 8'hFE; 14'h182D: rddata <= 8'h75; 14'h182E: rddata <= 8'h7E; 14'h182F: rddata <= 8'h18;
            14'h1830: rddata <= 8'h72; 14'h1831: rddata <= 8'h31; 14'h1832: rddata <= 8'h80; 14'h1833: rddata <= 8'h00;
            14'h1834: rddata <= 8'h00; 14'h1835: rddata <= 8'h00; 14'h1836: rddata <= 8'h81; 14'h1837: rddata <= 8'hCD;
            14'h1838: rddata <= 8'h13; 14'h1839: rddata <= 8'h15; 14'h183A: rddata <= 8'h11; 14'h183B: rddata <= 8'hC9;
            14'h183C: rddata <= 8'h13; 14'h183D: rddata <= 8'hD5; 14'h183E: rddata <= 8'hE5; 14'h183F: rddata <= 8'hCD;
            14'h1840: rddata <= 8'h2E; 14'h1841: rddata <= 8'h15; 14'h1842: rddata <= 8'hCD; 14'h1843: rddata <= 8'hCB;
            14'h1844: rddata <= 8'h13; 14'h1845: rddata <= 8'hE1; 14'h1846: rddata <= 8'hCD; 14'h1847: rddata <= 8'h13;
            14'h1848: rddata <= 8'h15; 14'h1849: rddata <= 8'h7E; 14'h184A: rddata <= 8'h23; 14'h184B: rddata <= 8'hCD;
            14'h184C: rddata <= 8'h20; 14'h184D: rddata <= 8'h15; 14'h184E: rddata <= 8'h06; 14'h184F: rddata <= 8'hF1;
            14'h1850: rddata <= 8'hC1; 14'h1851: rddata <= 8'hD1; 14'h1852: rddata <= 8'h3D; 14'h1853: rddata <= 8'hC8;
            14'h1854: rddata <= 8'hD5; 14'h1855: rddata <= 8'hC5; 14'h1856: rddata <= 8'hF5; 14'h1857: rddata <= 8'hE5;
            14'h1858: rddata <= 8'hCD; 14'h1859: rddata <= 8'hCB; 14'h185A: rddata <= 8'h13; 14'h185B: rddata <= 8'hE1;
            14'h185C: rddata <= 8'hCD; 14'h185D: rddata <= 8'h31; 14'h185E: rddata <= 8'h15; 14'h185F: rddata <= 8'hE5;
            14'h1860: rddata <= 8'hCD; 14'h1861: rddata <= 8'h61; 14'h1862: rddata <= 8'h12; 14'h1863: rddata <= 8'hE1;
            14'h1864: rddata <= 8'h18; 14'h1865: rddata <= 8'hE9; 14'h1866: rddata <= 8'hEF; 14'h1867: rddata <= 8'h21;
            14'h1868: rddata <= 8'h20; 14'h1869: rddata <= 8'h38; 14'h186A: rddata <= 8'hFA; 14'h186B: rddata <= 8'hC4;
            14'h186C: rddata <= 8'h18; 14'h186D: rddata <= 8'h21; 14'h186E: rddata <= 8'h41; 14'h186F: rddata <= 8'h38;
            14'h1870: rddata <= 8'hCD; 14'h1871: rddata <= 8'h20; 14'h1872: rddata <= 8'h15; 14'h1873: rddata <= 8'h21;
            14'h1874: rddata <= 8'h20; 14'h1875: rddata <= 8'h38; 14'h1876: rddata <= 8'hC8; 14'h1877: rddata <= 8'h86;
            14'h1878: rddata <= 8'hE6; 14'h1879: rddata <= 8'h07; 14'h187A: rddata <= 8'h06; 14'h187B: rddata <= 8'h00;
            14'h187C: rddata <= 8'h77; 14'h187D: rddata <= 8'h23; 14'h187E: rddata <= 8'h87; 14'h187F: rddata <= 8'h87;
            14'h1880: rddata <= 8'h4F; 14'h1881: rddata <= 8'h09; 14'h1882: rddata <= 8'hCD; 14'h1883: rddata <= 8'h31;
            14'h1884: rddata <= 8'h15; 14'h1885: rddata <= 8'hCD; 14'h1886: rddata <= 8'hCB; 14'h1887: rddata <= 8'h13;
            14'h1888: rddata <= 8'h3A; 14'h1889: rddata <= 8'h1F; 14'h188A: rddata <= 8'h38; 14'h188B: rddata <= 8'h3C;
            14'h188C: rddata <= 8'hE6; 14'h188D: rddata <= 8'h03; 14'h188E: rddata <= 8'h06; 14'h188F: rddata <= 8'h00;
            14'h1890: rddata <= 8'hFE; 14'h1891: rddata <= 8'h01; 14'h1892: rddata <= 8'h88; 14'h1893: rddata <= 8'h32;
            14'h1894: rddata <= 8'h1F; 14'h1895: rddata <= 8'h38; 14'h1896: rddata <= 8'h21; 14'h1897: rddata <= 8'hC7;
            14'h1898: rddata <= 8'h18; 14'h1899: rddata <= 8'h87; 14'h189A: rddata <= 8'h87; 14'h189B: rddata <= 8'h4F;
            14'h189C: rddata <= 8'h09; 14'h189D: rddata <= 8'hCD; 14'h189E: rddata <= 8'h53; 14'h189F: rddata <= 8'h12;
            14'h18A0: rddata <= 8'hCD; 14'h18A1: rddata <= 8'h2E; 14'h18A2: rddata <= 8'h15; 14'h18A3: rddata <= 8'h7B;
            14'h18A4: rddata <= 8'h59; 14'h18A5: rddata <= 8'hEE; 14'h18A6: rddata <= 8'h4F; 14'h18A7: rddata <= 8'h4F;
            14'h18A8: rddata <= 8'h36; 14'h18A9: rddata <= 8'h80; 14'h18AA: rddata <= 8'h2B; 14'h18AB: rddata <= 8'h46;
            14'h18AC: rddata <= 8'h36; 14'h18AD: rddata <= 8'h80; 14'h18AE: rddata <= 8'h21; 14'h18AF: rddata <= 8'h1E;
            14'h18B0: rddata <= 8'h38; 14'h18B1: rddata <= 8'h34; 14'h18B2: rddata <= 8'h7E; 14'h18B3: rddata <= 8'hD6;
            14'h18B4: rddata <= 8'hAB; 14'h18B5: rddata <= 8'h20; 14'h18B6: rddata <= 8'h04; 14'h18B7: rddata <= 8'h77;
            14'h18B8: rddata <= 8'h0C; 14'h18B9: rddata <= 8'h15; 14'h18BA: rddata <= 8'h1C; 14'h18BB: rddata <= 8'hCD;
            14'h18BC: rddata <= 8'hB0; 14'h18BD: rddata <= 8'h12; 14'h18BE: rddata <= 8'h21; 14'h18BF: rddata <= 8'h41;
            14'h18C0: rddata <= 8'h38; 14'h18C1: rddata <= 8'hC3; 14'h18C2: rddata <= 8'h3A; 14'h18C3: rddata <= 8'h15;
            14'h18C4: rddata <= 8'h77; 14'h18C5: rddata <= 8'h2B; 14'h18C6: rddata <= 8'h77; 14'h18C7: rddata <= 8'h2B;
            14'h18C8: rddata <= 8'h77; 14'h18C9: rddata <= 8'h18; 14'h18CA: rddata <= 8'hD5; 14'h18CB: rddata <= 8'h68;
            14'h18CC: rddata <= 8'hB1; 14'h18CD: rddata <= 8'h46; 14'h18CE: rddata <= 8'h68; 14'h18CF: rddata <= 8'h99;
            14'h18D0: rddata <= 8'hE9; 14'h18D1: rddata <= 8'h92; 14'h18D2: rddata <= 8'h69; 14'h18D3: rddata <= 8'h10;
            14'h18D4: rddata <= 8'hD1; 14'h18D5: rddata <= 8'h75; 14'h18D6: rddata <= 8'h68; 14'h18D7: rddata <= 8'h21;
            14'h18D8: rddata <= 8'h53; 14'h18D9: rddata <= 8'h19; 14'h18DA: rddata <= 8'hCD; 14'h18DB: rddata <= 8'h53;
            14'h18DC: rddata <= 8'h12; 14'h18DD: rddata <= 8'h3A; 14'h18DE: rddata <= 8'hE7; 14'h18DF: rddata <= 8'h38;
            14'h18E0: rddata <= 8'hFE; 14'h18E1: rddata <= 8'h77; 14'h18E2: rddata <= 8'hD8; 14'h18E3: rddata <= 8'h3A;
            14'h18E4: rddata <= 8'hE6; 14'h18E5: rddata <= 8'h38; 14'h18E6: rddata <= 8'hB7; 14'h18E7: rddata <= 8'hF2;
            14'h18E8: rddata <= 8'hF3; 14'h18E9: rddata <= 8'h18; 14'h18EA: rddata <= 8'hE6; 14'h18EB: rddata <= 8'h7F;
            14'h18EC: rddata <= 8'h32; 14'h18ED: rddata <= 8'hE6; 14'h18EE: rddata <= 8'h38; 14'h18EF: rddata <= 8'h11;
            14'h18F0: rddata <= 8'h0B; 14'h18F1: rddata <= 8'h15; 14'h18F2: rddata <= 8'hD5; 14'h18F3: rddata <= 8'h01;
            14'h18F4: rddata <= 8'h22; 14'h18F5: rddata <= 8'h7E; 14'h18F6: rddata <= 8'h11; 14'h18F7: rddata <= 8'h83;
            14'h18F8: rddata <= 8'hF9; 14'h18F9: rddata <= 8'hCD; 14'h18FA: rddata <= 8'hCB; 14'h18FB: rddata <= 8'h13;
            14'h18FC: rddata <= 8'hCD; 14'h18FD: rddata <= 8'h13; 14'h18FE: rddata <= 8'h15; 14'h18FF: rddata <= 8'hCD;
            14'h1900: rddata <= 8'hB1; 14'h1901: rddata <= 8'h15; 14'h1902: rddata <= 8'hC1; 14'h1903: rddata <= 8'hD1;
            14'h1904: rddata <= 8'hCD; 14'h1905: rddata <= 8'h5E; 14'h1906: rddata <= 8'h12; 14'h1907: rddata <= 8'h01;
            14'h1908: rddata <= 8'h00; 14'h1909: rddata <= 8'h7F; 14'h190A: rddata <= 8'h11; 14'h190B: rddata <= 8'h00;
            14'h190C: rddata <= 8'h00; 14'h190D: rddata <= 8'hCD; 14'h190E: rddata <= 8'h5B; 14'h190F: rddata <= 8'h15;
            14'h1910: rddata <= 8'hFA; 14'h1911: rddata <= 8'h35; 14'h1912: rddata <= 8'h19; 14'h1913: rddata <= 8'h01;
            14'h1914: rddata <= 8'h80; 14'h1915: rddata <= 8'h7F; 14'h1916: rddata <= 8'h11; 14'h1917: rddata <= 8'h00;
            14'h1918: rddata <= 8'h00; 14'h1919: rddata <= 8'hCD; 14'h191A: rddata <= 8'h61; 14'h191B: rddata <= 8'h12;
            14'h191C: rddata <= 8'h01; 14'h191D: rddata <= 8'h80; 14'h191E: rddata <= 8'h80; 14'h191F: rddata <= 8'h11;
            14'h1920: rddata <= 8'h00; 14'h1921: rddata <= 8'h00; 14'h1922: rddata <= 8'hCD; 14'h1923: rddata <= 8'h61;
            14'h1924: rddata <= 8'h12; 14'h1925: rddata <= 8'hEF; 14'h1926: rddata <= 8'hF4; 14'h1927: rddata <= 8'h0B;
            14'h1928: rddata <= 8'h15; 14'h1929: rddata <= 8'h01; 14'h192A: rddata <= 8'h00; 14'h192B: rddata <= 8'h7F;
            14'h192C: rddata <= 8'h11; 14'h192D: rddata <= 8'h00; 14'h192E: rddata <= 8'h00; 14'h192F: rddata <= 8'hCD;
            14'h1930: rddata <= 8'h61; 14'h1931: rddata <= 8'h12; 14'h1932: rddata <= 8'hCD; 14'h1933: rddata <= 8'h0B;
            14'h1934: rddata <= 8'h15; 14'h1935: rddata <= 8'h3A; 14'h1936: rddata <= 8'hE6; 14'h1937: rddata <= 8'h38;
            14'h1938: rddata <= 8'hB7; 14'h1939: rddata <= 8'hF5; 14'h193A: rddata <= 8'hF2; 14'h193B: rddata <= 8'h42;
            14'h193C: rddata <= 8'h19; 14'h193D: rddata <= 8'hEE; 14'h193E: rddata <= 8'h80; 14'h193F: rddata <= 8'h32;
            14'h1940: rddata <= 8'hE6; 14'h1941: rddata <= 8'h38; 14'h1942: rddata <= 8'h21; 14'h1943: rddata <= 8'h5B;
            14'h1944: rddata <= 8'h19; 14'h1945: rddata <= 8'hCD; 14'h1946: rddata <= 8'h37; 14'h1947: rddata <= 8'h18;
            14'h1948: rddata <= 8'hF1; 14'h1949: rddata <= 8'hF0; 14'h194A: rddata <= 8'h3A; 14'h194B: rddata <= 8'hE6;
            14'h194C: rddata <= 8'h38; 14'h194D: rddata <= 8'hEE; 14'h194E: rddata <= 8'h80; 14'h194F: rddata <= 8'h32;
            14'h1950: rddata <= 8'hE6; 14'h1951: rddata <= 8'h38; 14'h1952: rddata <= 8'hC9; 14'h1953: rddata <= 8'hDB;
            14'h1954: rddata <= 8'h0F; 14'h1955: rddata <= 8'h49; 14'h1956: rddata <= 8'h81; 14'h1957: rddata <= 8'h00;
            14'h1958: rddata <= 8'h00; 14'h1959: rddata <= 8'h00; 14'h195A: rddata <= 8'h7F; 14'h195B: rddata <= 8'h05;
            14'h195C: rddata <= 8'hFB; 14'h195D: rddata <= 8'hD7; 14'h195E: rddata <= 8'h1E; 14'h195F: rddata <= 8'h86;
            14'h1960: rddata <= 8'h65; 14'h1961: rddata <= 8'h26; 14'h1962: rddata <= 8'h99; 14'h1963: rddata <= 8'h87;
            14'h1964: rddata <= 8'h58; 14'h1965: rddata <= 8'h34; 14'h1966: rddata <= 8'h23; 14'h1967: rddata <= 8'h87;
            14'h1968: rddata <= 8'hE1; 14'h1969: rddata <= 8'h5D; 14'h196A: rddata <= 8'hA5; 14'h196B: rddata <= 8'h86;
            14'h196C: rddata <= 8'hDB; 14'h196D: rddata <= 8'h0F; 14'h196E: rddata <= 8'h49; 14'h196F: rddata <= 8'h83;
            14'h1970: rddata <= 8'hCD; 14'h1971: rddata <= 8'h13; 14'h1972: rddata <= 8'h15; 14'h1973: rddata <= 8'hCD;
            14'h1974: rddata <= 8'hDD; 14'h1975: rddata <= 8'h18; 14'h1976: rddata <= 8'hC1; 14'h1977: rddata <= 8'hE1;
            14'h1978: rddata <= 8'hCD; 14'h1979: rddata <= 8'h13; 14'h197A: rddata <= 8'h15; 14'h197B: rddata <= 8'hEB;
            14'h197C: rddata <= 8'hCD; 14'h197D: rddata <= 8'h23; 14'h197E: rddata <= 8'h15; 14'h197F: rddata <= 8'hCD;
            14'h1980: rddata <= 8'hD7; 14'h1981: rddata <= 8'h18; 14'h1982: rddata <= 8'hC3; 14'h1983: rddata <= 8'h2D;
            14'h1984: rddata <= 8'h14; 14'h1985: rddata <= 8'hF7; 14'h1986: rddata <= 8'h0E; 14'h1987: rddata <= 8'hC3;
            14'h1988: rddata <= 8'hC4; 14'h1989: rddata <= 8'h03; 14'h198A: rddata <= 8'hF7; 14'h198B: rddata <= 8'h0D;
            14'h198C: rddata <= 8'hF5; 14'h198D: rddata <= 8'h3A; 14'h198E: rddata <= 8'h47; 14'h198F: rddata <= 8'h38;
            14'h1990: rddata <= 8'hB7; 14'h1991: rddata <= 8'hCA; 14'h1992: rddata <= 8'hD6; 14'h1993: rddata <= 8'h19;
            14'h1994: rddata <= 8'hF1; 14'h1995: rddata <= 8'hF5; 14'h1996: rddata <= 8'hFE; 14'h1997: rddata <= 8'h09;
            14'h1998: rddata <= 8'h20; 14'h1999: rddata <= 8'h0C; 14'h199A: rddata <= 8'h3E; 14'h199B: rddata <= 8'h20;
            14'h199C: rddata <= 8'hDF; 14'h199D: rddata <= 8'h3A; 14'h199E: rddata <= 8'h46; 14'h199F: rddata <= 8'h38;
            14'h19A0: rddata <= 8'hE6; 14'h19A1: rddata <= 8'h07; 14'h19A2: rddata <= 8'h20; 14'h19A3: rddata <= 8'hF6;
            14'h19A4: rddata <= 8'hF1; 14'h19A5: rddata <= 8'hC9; 14'h19A6: rddata <= 8'hF1; 14'h19A7: rddata <= 8'hF5;
            14'h19A8: rddata <= 8'hD6; 14'h19A9: rddata <= 8'h0D; 14'h19AA: rddata <= 8'h28; 14'h19AB: rddata <= 8'h0B;
            14'h19AC: rddata <= 8'h38; 14'h19AD: rddata <= 8'h0C; 14'h19AE: rddata <= 8'h3A; 14'h19AF: rddata <= 8'h46;
            14'h19B0: rddata <= 8'h38; 14'h19B1: rddata <= 8'h3C; 14'h19B2: rddata <= 8'hFE; 14'h19B3: rddata <= 8'h84;
            14'h19B4: rddata <= 8'hCC; 14'h19B5: rddata <= 8'hC7; 14'h19B6: rddata <= 8'h19; 14'h19B7: rddata <= 8'h32;
            14'h19B8: rddata <= 8'h46; 14'h19B9: rddata <= 8'h38; 14'h19BA: rddata <= 8'hF1; 14'h19BB: rddata <= 8'hC3;
            14'h19BC: rddata <= 8'hE8; 14'h19BD: rddata <= 8'h1A; 14'h19BE: rddata <= 8'hAF; 14'h19BF: rddata <= 8'h32;
            14'h19C0: rddata <= 8'h47; 14'h19C1: rddata <= 8'h38; 14'h19C2: rddata <= 8'h3A; 14'h19C3: rddata <= 8'h46;
            14'h19C4: rddata <= 8'h38; 14'h19C5: rddata <= 8'hB7; 14'h19C6: rddata <= 8'hC8; 14'h19C7: rddata <= 8'h3E;
            14'h19C8: rddata <= 8'h0D; 14'h19C9: rddata <= 8'hCD; 14'h19CA: rddata <= 8'hBB; 14'h19CB: rddata <= 8'h19;
            14'h19CC: rddata <= 8'h3E; 14'h19CD: rddata <= 8'h0A; 14'h19CE: rddata <= 8'hCD; 14'h19CF: rddata <= 8'hBB;
            14'h19D0: rddata <= 8'h19; 14'h19D1: rddata <= 8'hAF; 14'h19D2: rddata <= 8'h32; 14'h19D3: rddata <= 8'h46;
            14'h19D4: rddata <= 8'h38; 14'h19D5: rddata <= 8'hC9; 14'h19D6: rddata <= 8'hF1; 14'h19D7: rddata <= 8'hC3;
            14'h19D8: rddata <= 8'h72; 14'h19D9: rddata <= 8'h1D; 14'h19DA: rddata <= 8'hCD; 14'h19DB: rddata <= 8'h2F;
            14'h19DC: rddata <= 8'h1A; 14'h19DD: rddata <= 8'hC9; 14'h19DE: rddata <= 8'h3A; 14'h19DF: rddata <= 8'h00;
            14'h19E0: rddata <= 8'h38; 14'h19E1: rddata <= 8'hB7; 14'h19E2: rddata <= 8'hC8; 14'h19E3: rddata <= 8'h18;
            14'h19E4: rddata <= 8'h05; 14'h19E5: rddata <= 8'h36; 14'h19E6: rddata <= 8'h00; 14'h19E7: rddata <= 8'h21;
            14'h19E8: rddata <= 8'h5F; 14'h19E9: rddata <= 8'h38; 14'h19EA: rddata <= 8'h3E; 14'h19EB: rddata <= 8'h0D;
            14'h19EC: rddata <= 8'hDF; 14'h19ED: rddata <= 8'h3E; 14'h19EE: rddata <= 8'h0A; 14'h19EF: rddata <= 8'hDF;
            14'h19F0: rddata <= 8'h3A; 14'h19F1: rddata <= 8'h47; 14'h19F2: rddata <= 8'h38; 14'h19F3: rddata <= 8'hB7;
            14'h19F4: rddata <= 8'h28; 14'h19F5: rddata <= 8'h04; 14'h19F6: rddata <= 8'hAF; 14'h19F7: rddata <= 8'h32;
            14'h19F8: rddata <= 8'h46; 14'h19F9: rddata <= 8'h38; 14'h19FA: rddata <= 8'hC9; 14'h19FB: rddata <= 8'hD7;
            14'h19FC: rddata <= 8'hE5; 14'h19FD: rddata <= 8'hCD; 14'h19FE: rddata <= 8'h18; 14'h19FF: rddata <= 8'h1A;
            14'h1A00: rddata <= 8'h28; 14'h1A01: rddata <= 8'h09; 14'h1A02: rddata <= 8'hF5; 14'h1A03: rddata <= 8'hCD;
            14'h1A04: rddata <= 8'h4E; 14'h1A05: rddata <= 8'h0E; 14'h1A06: rddata <= 8'hF1; 14'h1A07: rddata <= 8'h5F;
            14'h1A08: rddata <= 8'hCD; 14'h1A09: rddata <= 8'h19; 14'h1A0A: rddata <= 8'h10; 14'h1A0B: rddata <= 8'h21;
            14'h1A0C: rddata <= 8'h6D; 14'h1A0D: rddata <= 8'h03; 14'h1A0E: rddata <= 8'h22; 14'h1A0F: rddata <= 8'hE4;
            14'h1A10: rddata <= 8'h38; 14'h1A11: rddata <= 8'h3E; 14'h1A12: rddata <= 8'h01; 14'h1A13: rddata <= 8'h32;
            14'h1A14: rddata <= 8'hAB; 14'h1A15: rddata <= 8'h38; 14'h1A16: rddata <= 8'hE1; 14'h1A17: rddata <= 8'hC9;
            14'h1A18: rddata <= 8'hE5; 14'h1A19: rddata <= 8'h21; 14'h1A1A: rddata <= 8'h0A; 14'h1A1B: rddata <= 8'h38;
            14'h1A1C: rddata <= 8'h7E; 14'h1A1D: rddata <= 8'h36; 14'h1A1E: rddata <= 8'h00; 14'h1A1F: rddata <= 8'hB7;
            14'h1A20: rddata <= 8'hCC; 14'h1A21: rddata <= 8'h39; 14'h1A22: rddata <= 8'h1A; 14'h1A23: rddata <= 8'hE1;
            14'h1A24: rddata <= 8'hC9; 14'h1A25: rddata <= 8'hCD; 14'h1A26: rddata <= 8'h39; 14'h1A27: rddata <= 8'h1A;
            14'h1A28: rddata <= 8'hC8; 14'h1A29: rddata <= 8'h32; 14'h1A2A: rddata <= 8'h0A; 14'h1A2B: rddata <= 8'h38;
            14'h1A2C: rddata <= 8'hFE; 14'h1A2D: rddata <= 8'h13; 14'h1A2E: rddata <= 8'hC0; 14'h1A2F: rddata <= 8'hAF;
            14'h1A30: rddata <= 8'h32; 14'h1A31: rddata <= 8'h0A; 14'h1A32: rddata <= 8'h38; 14'h1A33: rddata <= 8'hCD;
            14'h1A34: rddata <= 8'h39; 14'h1A35: rddata <= 8'h1A; 14'h1A36: rddata <= 8'h28; 14'h1A37: rddata <= 8'hFB;
            14'h1A38: rddata <= 8'hC9; 14'h1A39: rddata <= 8'hCD; 14'h1A3A: rddata <= 8'h7E; 14'h1A3B: rddata <= 8'h1E;
            14'h1A3C: rddata <= 8'hFE; 14'h1A3D: rddata <= 8'h03; 14'h1A3E: rddata <= 8'h20; 14'h1A3F: rddata <= 8'h0A;
            14'h1A40: rddata <= 8'h3A; 14'h1A41: rddata <= 8'h5E; 14'h1A42: rddata <= 8'h38; 14'h1A43: rddata <= 8'hB7;
            14'h1A44: rddata <= 8'hCC; 14'h1A45: rddata <= 8'hBE; 14'h1A46: rddata <= 8'h0B; 14'h1A47: rddata <= 8'hC3;
            14'h1A48: rddata <= 8'hCE; 14'h1A49: rddata <= 8'h1F; 14'h1A4A: rddata <= 8'hB7; 14'h1A4B: rddata <= 8'hC9;
            14'h1A4C: rddata <= 8'hAF; 14'h1A4D: rddata <= 8'h18; 14'h1A4E: rddata <= 8'h02; 14'h1A4F: rddata <= 8'h3E;
            14'h1A50: rddata <= 8'h01; 14'h1A51: rddata <= 8'h08; 14'h1A52: rddata <= 8'hCD; 14'h1A53: rddata <= 8'h7F;
            14'h1A54: rddata <= 8'h1A; 14'h1A55: rddata <= 8'hCD; 14'h1A56: rddata <= 8'h8E; 14'h1A57: rddata <= 8'h1A;
            14'h1A58: rddata <= 8'h28; 14'h1A59: rddata <= 8'h02; 14'h1A5A: rddata <= 8'h36; 14'h1A5B: rddata <= 8'hA0;
            14'h1A5C: rddata <= 8'h08; 14'h1A5D: rddata <= 8'hB7; 14'h1A5E: rddata <= 8'h1A; 14'h1A5F: rddata <= 8'h20;
            14'h1A60: rddata <= 8'h03; 14'h1A61: rddata <= 8'h2F; 14'h1A62: rddata <= 8'hA6; 14'h1A63: rddata <= 8'h06;
            14'h1A64: rddata <= 8'hB6; 14'h1A65: rddata <= 8'h77; 14'h1A66: rddata <= 8'hE1; 14'h1A67: rddata <= 8'hC9;
            14'h1A68: rddata <= 8'hD7; 14'h1A69: rddata <= 8'hCD; 14'h1A6A: rddata <= 8'h7F; 14'h1A6B: rddata <= 8'h1A;
            14'h1A6C: rddata <= 8'hCD; 14'h1A6D: rddata <= 8'h8E; 14'h1A6E: rddata <= 8'h1A; 14'h1A6F: rddata <= 8'h20;
            14'h1A70: rddata <= 8'h06; 14'h1A71: rddata <= 8'h1A; 14'h1A72: rddata <= 8'hA6; 14'h1A73: rddata <= 8'h16;
            14'h1A74: rddata <= 8'h01; 14'h1A75: rddata <= 8'h20; 14'h1A76: rddata <= 8'h02; 14'h1A77: rddata <= 8'h16;
            14'h1A78: rddata <= 8'h00; 14'h1A79: rddata <= 8'hAF; 14'h1A7A: rddata <= 8'hCD; 14'h1A7B: rddata <= 8'h23;
            14'h1A7C: rddata <= 8'h0B; 14'h1A7D: rddata <= 8'hE1; 14'h1A7E: rddata <= 8'hC9; 14'h1A7F: rddata <= 8'hCF;
            14'h1A80: rddata <= 8'h28; 14'h1A81: rddata <= 8'hCD; 14'h1A82: rddata <= 8'hD0; 14'h1A83: rddata <= 8'h1A;
            14'h1A84: rddata <= 8'hD5; 14'h1A85: rddata <= 8'hCF; 14'h1A86: rddata <= 8'h2C; 14'h1A87: rddata <= 8'hCD;
            14'h1A88: rddata <= 8'hD0; 14'h1A89: rddata <= 8'h1A; 14'h1A8A: rddata <= 8'hCF; 14'h1A8B: rddata <= 8'h29;
            14'h1A8C: rddata <= 8'hC1; 14'h1A8D: rddata <= 8'hC9; 14'h1A8E: rddata <= 8'hE3; 14'h1A8F: rddata <= 8'hE5;
            14'h1A90: rddata <= 8'hC5; 14'h1A91: rddata <= 8'hD5; 14'h1A92: rddata <= 8'h21; 14'h1A93: rddata <= 8'h47;
            14'h1A94: rddata <= 8'h00; 14'h1A95: rddata <= 8'hE7; 14'h1A96: rddata <= 8'hDA; 14'h1A97: rddata <= 8'h97;
            14'h1A98: rddata <= 8'h06; 14'h1A99: rddata <= 8'h21; 14'h1A9A: rddata <= 8'h4F; 14'h1A9B: rddata <= 8'h00;
            14'h1A9C: rddata <= 8'hC5; 14'h1A9D: rddata <= 8'hD1; 14'h1A9E: rddata <= 8'hE7; 14'h1A9F: rddata <= 8'h38;
            14'h1AA0: rddata <= 8'hF5; 14'h1AA1: rddata <= 8'hD1; 14'h1AA2: rddata <= 8'hC1; 14'h1AA3: rddata <= 8'h21;
            14'h1AA4: rddata <= 8'h28; 14'h1AA5: rddata <= 8'h30; 14'h1AA6: rddata <= 8'h7B; 14'h1AA7: rddata <= 8'h11;
            14'h1AA8: rddata <= 8'h28; 14'h1AA9: rddata <= 8'h00; 14'h1AAA: rddata <= 8'hFE; 14'h1AAB: rddata <= 8'h03;
            14'h1AAC: rddata <= 8'h38; 14'h1AAD: rddata <= 8'h06; 14'h1AAE: rddata <= 8'h19; 14'h1AAF: rddata <= 8'h3D;
            14'h1AB0: rddata <= 8'h3D; 14'h1AB1: rddata <= 8'h3D; 14'h1AB2: rddata <= 8'h18; 14'h1AB3: rddata <= 8'hF6;
            14'h1AB4: rddata <= 8'h07; 14'h1AB5: rddata <= 8'hCB; 14'h1AB6: rddata <= 8'h29; 14'h1AB7: rddata <= 8'h30;
            14'h1AB8: rddata <= 8'h01; 14'h1AB9: rddata <= 8'h3C; 14'h1ABA: rddata <= 8'h09; 14'h1ABB: rddata <= 8'h11;
            14'h1ABC: rddata <= 8'hCA; 14'h1ABD: rddata <= 8'h1A; 14'h1ABE: rddata <= 8'hB7; 14'h1ABF: rddata <= 8'h28;
            14'h1AC0: rddata <= 8'h04; 14'h1AC1: rddata <= 8'h13; 14'h1AC2: rddata <= 8'h3D; 14'h1AC3: rddata <= 8'h18;
            14'h1AC4: rddata <= 8'hF9; 14'h1AC5: rddata <= 8'h7E; 14'h1AC6: rddata <= 8'hF6; 14'h1AC7: rddata <= 8'hA0;
            14'h1AC8: rddata <= 8'hAE; 14'h1AC9: rddata <= 8'hC9; 14'h1ACA: rddata <= 8'h01; 14'h1ACB: rddata <= 8'h02;
            14'h1ACC: rddata <= 8'h04; 14'h1ACD: rddata <= 8'h08; 14'h1ACE: rddata <= 8'h10; 14'h1ACF: rddata <= 8'h40;
            14'h1AD0: rddata <= 8'hCD; 14'h1AD1: rddata <= 8'h85; 14'h1AD2: rddata <= 8'h09; 14'h1AD3: rddata <= 8'hC3;
            14'h1AD4: rddata <= 8'h82; 14'h1AD5: rddata <= 8'h06; 14'h1AD6: rddata <= 8'hD5; 14'h1AD7: rddata <= 8'hCD;
            14'h1AD8: rddata <= 8'h7F; 14'h1AD9: rddata <= 8'h1A; 14'h1ADA: rddata <= 8'hE5; 14'h1ADB: rddata <= 8'hCD;
            14'h1ADC: rddata <= 8'h64; 14'h1ADD: rddata <= 8'h1E; 14'h1ADE: rddata <= 8'hE1; 14'h1ADF: rddata <= 8'hD1;
            14'h1AE0: rddata <= 8'hC9; 14'h1AE1: rddata <= 8'h3E; 14'h1AE2: rddata <= 8'h0D; 14'h1AE3: rddata <= 8'hCD;
            14'h1AE4: rddata <= 8'hE8; 14'h1AE5: rddata <= 8'h1A; 14'h1AE6: rddata <= 8'h3E; 14'h1AE7: rddata <= 8'h0A;
            14'h1AE8: rddata <= 8'hF7; 14'h1AE9: rddata <= 8'h11; 14'h1AEA: rddata <= 8'hF5; 14'h1AEB: rddata <= 8'hF5;
            14'h1AEC: rddata <= 8'hD9; 14'h1AED: rddata <= 8'hDB; 14'h1AEE: rddata <= 8'hFE; 14'h1AEF: rddata <= 8'hE6;
            14'h1AF0: rddata <= 8'h01; 14'h1AF1: rddata <= 8'h28; 14'h1AF2: rddata <= 8'hFA; 14'h1AF3: rddata <= 8'hCD;
            14'h1AF4: rddata <= 8'h08; 14'h1AF5: rddata <= 8'h1B; 14'h1AF6: rddata <= 8'h1E; 14'h1AF7: rddata <= 8'h08;
            14'h1AF8: rddata <= 8'hF1; 14'h1AF9: rddata <= 8'hCD; 14'h1AFA: rddata <= 8'h0A; 14'h1AFB: rddata <= 8'h1B;
            14'h1AFC: rddata <= 8'h0F; 14'h1AFD: rddata <= 8'h1D; 14'h1AFE: rddata <= 8'h20; 14'h1AFF: rddata <= 8'hF9;
            14'h1B00: rddata <= 8'h3E; 14'h1B01: rddata <= 8'h01; 14'h1B02: rddata <= 8'hCD; 14'h1B03: rddata <= 8'h0A;
            14'h1B04: rddata <= 8'h1B; 14'h1B05: rddata <= 8'hD9; 14'h1B06: rddata <= 8'hF1; 14'h1B07: rddata <= 8'hC9;
            14'h1B08: rddata <= 8'h3E; 14'h1B09: rddata <= 8'h00; 14'h1B0A: rddata <= 8'hD3; 14'h1B0B: rddata <= 8'hFE;
            14'h1B0C: rddata <= 8'h26; 14'h1B0D: rddata <= 8'hB1; 14'h1B0E: rddata <= 8'h25; 14'h1B0F: rddata <= 8'h20;
            14'h1B10: rddata <= 8'hFD; 14'h1B11: rddata <= 8'h00; 14'h1B12: rddata <= 8'h00; 14'h1B13: rddata <= 8'h00;
            14'h1B14: rddata <= 8'hC9; 14'h1B15: rddata <= 8'hE5; 14'h1B16: rddata <= 8'hD5; 14'h1B17: rddata <= 8'hCD;
            14'h1B18: rddata <= 8'hE1; 14'h1B19: rddata <= 8'h1A; 14'h1B1A: rddata <= 8'h21; 14'h1B1B: rddata <= 8'h28;
            14'h1B1C: rddata <= 8'h30; 14'h1B1D: rddata <= 8'h11; 14'h1B1E: rddata <= 8'hE8; 14'h1B1F: rddata <= 8'h33;
            14'h1B20: rddata <= 8'h7E; 14'h1B21: rddata <= 8'hCD; 14'h1B22: rddata <= 8'hE8; 14'h1B23: rddata <= 8'h1A;
            14'h1B24: rddata <= 8'h23; 14'h1B25: rddata <= 8'hE7; 14'h1B26: rddata <= 8'h38; 14'h1B27: rddata <= 8'hF8;
            14'h1B28: rddata <= 8'hCD; 14'h1B29: rddata <= 8'hE1; 14'h1B2A: rddata <= 8'h1A; 14'h1B2B: rddata <= 8'hD1;
            14'h1B2C: rddata <= 8'hE1; 14'h1B2D: rddata <= 8'hC9; 14'h1B2E: rddata <= 8'hE5; 14'h1B2F: rddata <= 8'hD5;
            14'h1B30: rddata <= 8'hC5; 14'h1B31: rddata <= 8'h21; 14'h1B32: rddata <= 8'hE8; 14'h1B33: rddata <= 8'h1B;
            14'h1B34: rddata <= 8'hF5; 14'h1B35: rddata <= 8'hCD; 14'h1B36: rddata <= 8'h9D; 14'h1B37: rddata <= 8'h0E;
            14'h1B38: rddata <= 8'h21; 14'h1B39: rddata <= 8'hB5; 14'h1B3A: rddata <= 8'h00; 14'h1B3B: rddata <= 8'hCD;
            14'h1B3C: rddata <= 8'h9D; 14'h1B3D: rddata <= 8'h0E; 14'h1B3E: rddata <= 8'hCD; 14'h1B3F: rddata <= 8'h7E;
            14'h1B40: rddata <= 8'h1E; 14'h1B41: rddata <= 8'hFE; 14'h1B42: rddata <= 8'h0D; 14'h1B43: rddata <= 8'h20;
            14'h1B44: rddata <= 8'hF9; 14'h1B45: rddata <= 8'hCD; 14'h1B46: rddata <= 8'hEA; 14'h1B47: rddata <= 8'h19;
            14'h1B48: rddata <= 8'hF1; 14'h1B49: rddata <= 8'hC1; 14'h1B4A: rddata <= 8'hD1; 14'h1B4B: rddata <= 8'hE1;
            14'h1B4C: rddata <= 8'hC9; 14'h1B4D: rddata <= 8'hD9; 14'h1B4E: rddata <= 8'h0E; 14'h1B4F: rddata <= 8'hFC;
            14'h1B50: rddata <= 8'hCD; 14'h1B51: rddata <= 8'h62; 14'h1B52: rddata <= 8'h1B; 14'h1B53: rddata <= 8'h38;
            14'h1B54: rddata <= 8'hFB; 14'h1B55: rddata <= 8'h26; 14'h1B56: rddata <= 8'h08; 14'h1B57: rddata <= 8'hCD;
            14'h1B58: rddata <= 8'h62; 14'h1B59: rddata <= 8'h1B; 14'h1B5A: rddata <= 8'hCB; 14'h1B5B: rddata <= 8'h15;
            14'h1B5C: rddata <= 8'h25; 14'h1B5D: rddata <= 8'h20; 14'h1B5E: rddata <= 8'hF8; 14'h1B5F: rddata <= 8'h7D;
            14'h1B60: rddata <= 8'hD9; 14'h1B61: rddata <= 8'hC9; 14'h1B62: rddata <= 8'hED; 14'h1B63: rddata <= 8'h78;
            14'h1B64: rddata <= 8'h1F; 14'h1B65: rddata <= 8'h38; 14'h1B66: rddata <= 8'hFB; 14'h1B67: rddata <= 8'hED;
            14'h1B68: rddata <= 8'h78; 14'h1B69: rddata <= 8'h1F; 14'h1B6A: rddata <= 8'h30; 14'h1B6B: rddata <= 8'hFB;
            14'h1B6C: rddata <= 8'hAF; 14'h1B6D: rddata <= 8'h3C; 14'h1B6E: rddata <= 8'hED; 14'h1B6F: rddata <= 8'h40;
            14'h1B70: rddata <= 8'hCB; 14'h1B71: rddata <= 8'h18; 14'h1B72: rddata <= 8'h38; 14'h1B73: rddata <= 8'hF9;
            14'h1B74: rddata <= 8'h3C; 14'h1B75: rddata <= 8'hED; 14'h1B76: rddata <= 8'h40; 14'h1B77: rddata <= 8'hCB;
            14'h1B78: rddata <= 8'h18; 14'h1B79: rddata <= 8'h30; 14'h1B7A: rddata <= 8'hF9; 14'h1B7B: rddata <= 8'hFE;
            14'h1B7C: rddata <= 8'h49; 14'h1B7D: rddata <= 8'hC9; 14'h1B7E: rddata <= 8'hC9; 14'h1B7F: rddata <= 8'hE5;
            14'h1B80: rddata <= 8'hD5; 14'h1B81: rddata <= 8'hC5; 14'h1B82: rddata <= 8'h21; 14'h1B83: rddata <= 8'hF7;
            14'h1B84: rddata <= 8'h1B; 14'h1B85: rddata <= 8'h18; 14'h1B86: rddata <= 8'hAD; 14'h1B87: rddata <= 8'hCD;
            14'h1B88: rddata <= 8'h8A; 14'h1B89: rddata <= 8'h1B; 14'h1B8A: rddata <= 8'hF5; 14'h1B8B: rddata <= 8'hD9;
            14'h1B8C: rddata <= 8'h0E; 14'h1B8D: rddata <= 8'hFC; 14'h1B8E: rddata <= 8'hF5; 14'h1B8F: rddata <= 8'hAF;
            14'h1B90: rddata <= 8'h1E; 14'h1B91: rddata <= 8'h01; 14'h1B92: rddata <= 8'hCD; 14'h1B93: rddata <= 8'hA5;
            14'h1B94: rddata <= 8'h1B; 14'h1B95: rddata <= 8'hF1; 14'h1B96: rddata <= 8'h1E; 14'h1B97: rddata <= 8'h08;
            14'h1B98: rddata <= 8'hCD; 14'h1B99: rddata <= 8'hA5; 14'h1B9A: rddata <= 8'h1B; 14'h1B9B: rddata <= 8'h3E;
            14'h1B9C: rddata <= 8'hFF; 14'h1B9D: rddata <= 8'h1E; 14'h1B9E: rddata <= 8'h02; 14'h1B9F: rddata <= 8'hCD;
            14'h1BA0: rddata <= 8'hA5; 14'h1BA1: rddata <= 8'h1B; 14'h1BA2: rddata <= 8'hD9; 14'h1BA3: rddata <= 8'hF1;
            14'h1BA4: rddata <= 8'hC9; 14'h1BA5: rddata <= 8'h17; 14'h1BA6: rddata <= 8'h2E; 14'h1BA7: rddata <= 8'h40;
            14'h1BA8: rddata <= 8'h38; 14'h1BA9: rddata <= 8'h02; 14'h1BAA: rddata <= 8'h2E; 14'h1BAB: rddata <= 8'h80;
            14'h1BAC: rddata <= 8'h06; 14'h1BAD: rddata <= 8'h04; 14'h1BAE: rddata <= 8'hED; 14'h1BAF: rddata <= 8'h41;
            14'h1BB0: rddata <= 8'h65; 14'h1BB1: rddata <= 8'h25; 14'h1BB2: rddata <= 8'h20; 14'h1BB3: rddata <= 8'hFD;
            14'h1BB4: rddata <= 8'h05; 14'h1BB5: rddata <= 8'h20; 14'h1BB6: rddata <= 8'hF7; 14'h1BB7: rddata <= 8'h1D;
            14'h1BB8: rddata <= 8'h20; 14'h1BB9: rddata <= 8'hEB; 14'h1BBA: rddata <= 8'hC9; 14'h1BBB: rddata <= 8'hC9;
            14'h1BBC: rddata <= 8'hF5; 14'h1BBD: rddata <= 8'hC5; 14'h1BBE: rddata <= 8'h06; 14'h1BBF: rddata <= 8'h0C;
            14'h1BC0: rddata <= 8'h3E; 14'h1BC1: rddata <= 8'hFF; 14'h1BC2: rddata <= 8'hCD; 14'h1BC3: rddata <= 8'h8A;
            14'h1BC4: rddata <= 8'h1B; 14'h1BC5: rddata <= 8'h10; 14'h1BC6: rddata <= 8'hF9; 14'h1BC7: rddata <= 8'hAF;
            14'h1BC8: rddata <= 8'hCD; 14'h1BC9: rddata <= 8'h8A; 14'h1BCA: rddata <= 8'h1B; 14'h1BCB: rddata <= 8'hC1;
            14'h1BCC: rddata <= 8'hF1; 14'h1BCD: rddata <= 8'hC9; 14'h1BCE: rddata <= 8'hF5; 14'h1BCF: rddata <= 8'hC5;
            14'h1BD0: rddata <= 8'h06; 14'h1BD1: rddata <= 8'h06; 14'h1BD2: rddata <= 8'hCD; 14'h1BD3: rddata <= 8'h4D;
            14'h1BD4: rddata <= 8'h1B; 14'h1BD5: rddata <= 8'h3C; 14'h1BD6: rddata <= 8'h20; 14'h1BD7: rddata <= 8'hF8;
            14'h1BD8: rddata <= 8'h10; 14'h1BD9: rddata <= 8'hF8; 14'h1BDA: rddata <= 8'hCD; 14'h1BDB: rddata <= 8'h4D;
            14'h1BDC: rddata <= 8'h1B; 14'h1BDD: rddata <= 8'hB7; 14'h1BDE: rddata <= 8'h28; 14'h1BDF: rddata <= 8'h05;
            14'h1BE0: rddata <= 8'h3C; 14'h1BE1: rddata <= 8'h28; 14'h1BE2: rddata <= 8'hF7; 14'h1BE3: rddata <= 8'h18;
            14'h1BE4: rddata <= 8'hEB; 14'h1BE5: rddata <= 8'hC1; 14'h1BE6: rddata <= 8'hF1; 14'h1BE7: rddata <= 8'hC9;
            14'h1BE8: rddata <= 8'h50; 14'h1BE9: rddata <= 8'h72; 14'h1BEA: rddata <= 8'h65; 14'h1BEB: rddata <= 8'h73;
            14'h1BEC: rddata <= 8'h73; 14'h1BED: rddata <= 8'h20; 14'h1BEE: rddata <= 8'h3C; 14'h1BEF: rddata <= 8'h50;
            14'h1BF0: rddata <= 8'h4C; 14'h1BF1: rddata <= 8'h41; 14'h1BF2: rddata <= 8'h59; 14'h1BF3: rddata <= 8'h3E;
            14'h1BF4: rddata <= 8'h0D; 14'h1BF5: rddata <= 8'h0A; 14'h1BF6: rddata <= 8'h00; 14'h1BF7: rddata <= 8'h50;
            14'h1BF8: rddata <= 8'h72; 14'h1BF9: rddata <= 8'h65; 14'h1BFA: rddata <= 8'h73; 14'h1BFB: rddata <= 8'h73;
            14'h1BFC: rddata <= 8'h20; 14'h1BFD: rddata <= 8'h3C; 14'h1BFE: rddata <= 8'h52; 14'h1BFF: rddata <= 8'h45;
            14'h1C00: rddata <= 8'h43; 14'h1C01: rddata <= 8'h4F; 14'h1C02: rddata <= 8'h52; 14'h1C03: rddata <= 8'h44;
            14'h1C04: rddata <= 8'h3E; 14'h1C05: rddata <= 8'h0D; 14'h1C06: rddata <= 8'h0A; 14'h1C07: rddata <= 8'h00;
            14'h1C08: rddata <= 8'hF7; 14'h1C09: rddata <= 8'h15; 14'h1C0A: rddata <= 8'hFE; 14'h1C0B: rddata <= 8'hAA;
            14'h1C0C: rddata <= 8'hCA; 14'h1C0D: rddata <= 8'h62; 14'h1C0E: rddata <= 8'h0C; 14'h1C0F: rddata <= 8'hCD;
            14'h1C10: rddata <= 8'hB8; 14'h1C11: rddata <= 8'h1C; 14'h1C12: rddata <= 8'hE5; 14'h1C13: rddata <= 8'hCD;
            14'h1C14: rddata <= 8'h25; 14'h1C15: rddata <= 8'h1D; 14'h1C16: rddata <= 8'h2A; 14'h1C17: rddata <= 8'h4F;
            14'h1C18: rddata <= 8'h38; 14'h1C19: rddata <= 8'hCD; 14'h1C1A: rddata <= 8'h38; 14'h1C1B: rddata <= 8'h1D;
            14'h1C1C: rddata <= 8'h06; 14'h1C1D: rddata <= 8'h0F; 14'h1C1E: rddata <= 8'hAF; 14'h1C1F: rddata <= 8'hCD;
            14'h1C20: rddata <= 8'h8A; 14'h1C21: rddata <= 8'h1B; 14'h1C22: rddata <= 8'h10; 14'h1C23: rddata <= 8'hFB;
            14'h1C24: rddata <= 8'h01; 14'h1C25: rddata <= 8'h40; 14'h1C26: rddata <= 8'h1F; 14'h1C27: rddata <= 8'hCD;
            14'h1C28: rddata <= 8'h4B; 14'h1C29: rddata <= 8'h1D; 14'h1C2A: rddata <= 8'hE1; 14'h1C2B: rddata <= 8'hC9;
            14'h1C2C: rddata <= 8'hF7; 14'h1C2D: rddata <= 8'h14; 14'h1C2E: rddata <= 8'hFE; 14'h1C2F: rddata <= 8'hAA;
            14'h1C30: rddata <= 8'hCA; 14'h1C31: rddata <= 8'h63; 14'h1C32: rddata <= 8'h0C; 14'h1C33: rddata <= 8'hD6;
            14'h1C34: rddata <= 8'h95; 14'h1C35: rddata <= 8'h28; 14'h1C36: rddata <= 8'h02; 14'h1C37: rddata <= 8'hAF;
            14'h1C38: rddata <= 8'h01; 14'h1C39: rddata <= 8'h2F; 14'h1C3A: rddata <= 8'h23; 14'h1C3B: rddata <= 8'hFE;
            14'h1C3C: rddata <= 8'h01; 14'h1C3D: rddata <= 8'hF5; 14'h1C3E: rddata <= 8'h3E; 14'h1C3F: rddata <= 8'hFF;
            14'h1C40: rddata <= 8'h32; 14'h1C41: rddata <= 8'h5E; 14'h1C42: rddata <= 8'h38; 14'h1C43: rddata <= 8'hCD;
            14'h1C44: rddata <= 8'hB1; 14'h1C45: rddata <= 8'h1C; 14'h1C46: rddata <= 8'hAF; 14'h1C47: rddata <= 8'h32;
            14'h1C48: rddata <= 8'h5D; 14'h1C49: rddata <= 8'h38; 14'h1C4A: rddata <= 8'hD5; 14'h1C4B: rddata <= 8'hCD;
            14'h1C4C: rddata <= 8'h2E; 14'h1C4D: rddata <= 8'h1B; 14'h1C4E: rddata <= 8'hCD; 14'h1C4F: rddata <= 8'hD9;
            14'h1C50: rddata <= 8'h1C; 14'h1C51: rddata <= 8'h21; 14'h1C52: rddata <= 8'h57; 14'h1C53: rddata <= 8'h38;
            14'h1C54: rddata <= 8'hCD; 14'h1C55: rddata <= 8'hED; 14'h1C56: rddata <= 8'h1C; 14'h1C57: rddata <= 8'hD1;
            14'h1C58: rddata <= 8'h28; 14'h1C59: rddata <= 8'h12; 14'h1C5A: rddata <= 8'h21; 14'h1C5B: rddata <= 8'h06;
            14'h1C5C: rddata <= 8'h1D; 14'h1C5D: rddata <= 8'hCD; 14'h1C5E: rddata <= 8'h0D; 14'h1C5F: rddata <= 8'h1D;
            14'h1C60: rddata <= 8'h06; 14'h1C61: rddata <= 8'h0A; 14'h1C62: rddata <= 8'hCD; 14'h1C63: rddata <= 8'h4D;
            14'h1C64: rddata <= 8'h1B; 14'h1C65: rddata <= 8'hB7; 14'h1C66: rddata <= 8'h20; 14'h1C67: rddata <= 8'hF8;
            14'h1C68: rddata <= 8'h10; 14'h1C69: rddata <= 8'hF8; 14'h1C6A: rddata <= 8'h18; 14'h1C6B: rddata <= 8'hDA;
            14'h1C6C: rddata <= 8'h21; 14'h1C6D: rddata <= 8'hFE; 14'h1C6E: rddata <= 8'h1C; 14'h1C6F: rddata <= 8'hCD;
            14'h1C70: rddata <= 8'h0D; 14'h1C71: rddata <= 8'h1D; 14'h1C72: rddata <= 8'hF1; 14'h1C73: rddata <= 8'h32;
            14'h1C74: rddata <= 8'hE4; 14'h1C75: rddata <= 8'h38; 14'h1C76: rddata <= 8'hDC; 14'h1C77: rddata <= 8'hBE;
            14'h1C78: rddata <= 8'h0B; 14'h1C79: rddata <= 8'h3A; 14'h1C7A: rddata <= 8'hE4; 14'h1C7B: rddata <= 8'h38;
            14'h1C7C: rddata <= 8'hFE; 14'h1C7D: rddata <= 8'h01; 14'h1C7E: rddata <= 8'h32; 14'h1C7F: rddata <= 8'h5E;
            14'h1C80: rddata <= 8'h38; 14'h1C81: rddata <= 8'h2A; 14'h1C82: rddata <= 8'h4F; 14'h1C83: rddata <= 8'h38;
            14'h1C84: rddata <= 8'hCD; 14'h1C85: rddata <= 8'h51; 14'h1C86: rddata <= 8'h1D; 14'h1C87: rddata <= 8'h20;
            14'h1C88: rddata <= 8'h11; 14'h1C89: rddata <= 8'h22; 14'h1C8A: rddata <= 8'hD6; 14'h1C8B: rddata <= 8'h38;
            14'h1C8C: rddata <= 8'h21; 14'h1C8D: rddata <= 8'h6E; 14'h1C8E: rddata <= 8'h03; 14'h1C8F: rddata <= 8'hCD;
            14'h1C90: rddata <= 8'h9D; 14'h1C91: rddata <= 8'h0E; 14'h1C92: rddata <= 8'h3E; 14'h1C93: rddata <= 8'hFF;
            14'h1C94: rddata <= 8'h32; 14'h1C95: rddata <= 8'h5E; 14'h1C96: rddata <= 8'h38; 14'h1C97: rddata <= 8'hC3;
            14'h1C98: rddata <= 8'h80; 14'h1C99: rddata <= 8'h04; 14'h1C9A: rddata <= 8'h23; 14'h1C9B: rddata <= 8'hEB;
            14'h1C9C: rddata <= 8'h2A; 14'h1C9D: rddata <= 8'hD6; 14'h1C9E: rddata <= 8'h38; 14'h1C9F: rddata <= 8'hE7;
            14'h1CA0: rddata <= 8'h38; 14'h1CA1: rddata <= 8'hEA; 14'h1CA2: rddata <= 8'h21; 14'h1CA3: rddata <= 8'hAB;
            14'h1CA4: rddata <= 8'h1C; 14'h1CA5: rddata <= 8'hCD; 14'h1CA6: rddata <= 8'h9D; 14'h1CA7: rddata <= 8'h0E;
            14'h1CA8: rddata <= 8'hC3; 14'h1CA9: rddata <= 8'h01; 14'h1CAA: rddata <= 8'h04; 14'h1CAB: rddata <= 8'h42;
            14'h1CAC: rddata <= 8'h61; 14'h1CAD: rddata <= 8'h64; 14'h1CAE: rddata <= 8'h0D; 14'h1CAF: rddata <= 8'h0A;
            14'h1CB0: rddata <= 8'h00; 14'h1CB1: rddata <= 8'hAF; 14'h1CB2: rddata <= 8'h32; 14'h1CB3: rddata <= 8'h51;
            14'h1CB4: rddata <= 8'h38; 14'h1CB5: rddata <= 8'h2B; 14'h1CB6: rddata <= 8'hD7; 14'h1CB7: rddata <= 8'hC8;
            14'h1CB8: rddata <= 8'hCD; 14'h1CB9: rddata <= 8'h85; 14'h1CBA: rddata <= 8'h09; 14'h1CBB: rddata <= 8'hE5;
            14'h1CBC: rddata <= 8'hCD; 14'h1CBD: rddata <= 8'h06; 14'h1CBE: rddata <= 8'h10; 14'h1CBF: rddata <= 8'h2B;
            14'h1CC0: rddata <= 8'h2B; 14'h1CC1: rddata <= 8'h2B; 14'h1CC2: rddata <= 8'h46; 14'h1CC3: rddata <= 8'h0E;
            14'h1CC4: rddata <= 8'h06; 14'h1CC5: rddata <= 8'h21; 14'h1CC6: rddata <= 8'h51; 14'h1CC7: rddata <= 8'h38;
            14'h1CC8: rddata <= 8'h1A; 14'h1CC9: rddata <= 8'h77; 14'h1CCA: rddata <= 8'h23; 14'h1CCB: rddata <= 8'h13;
            14'h1CCC: rddata <= 8'h0D; 14'h1CCD: rddata <= 8'h28; 14'h1CCE: rddata <= 8'h08; 14'h1CCF: rddata <= 8'h10;
            14'h1CD0: rddata <= 8'hF7; 14'h1CD1: rddata <= 8'h41; 14'h1CD2: rddata <= 8'h36; 14'h1CD3: rddata <= 8'h00;
            14'h1CD4: rddata <= 8'h23; 14'h1CD5: rddata <= 8'h10; 14'h1CD6: rddata <= 8'hFB; 14'h1CD7: rddata <= 8'hE1;
            14'h1CD8: rddata <= 8'hC9; 14'h1CD9: rddata <= 8'hCD; 14'h1CDA: rddata <= 8'hCE; 14'h1CDB: rddata <= 8'h1B;
            14'h1CDC: rddata <= 8'hAF; 14'h1CDD: rddata <= 8'h32; 14'h1CDE: rddata <= 8'h5D; 14'h1CDF: rddata <= 8'h38;
            14'h1CE0: rddata <= 8'h21; 14'h1CE1: rddata <= 8'h57; 14'h1CE2: rddata <= 8'h38; 14'h1CE3: rddata <= 8'h06;
            14'h1CE4: rddata <= 8'h06; 14'h1CE5: rddata <= 8'hCD; 14'h1CE6: rddata <= 8'h4D; 14'h1CE7: rddata <= 8'h1B;
            14'h1CE8: rddata <= 8'h77; 14'h1CE9: rddata <= 8'h23; 14'h1CEA: rddata <= 8'h10; 14'h1CEB: rddata <= 8'hF9;
            14'h1CEC: rddata <= 8'hC9; 14'h1CED: rddata <= 8'h01; 14'h1CEE: rddata <= 8'h51; 14'h1CEF: rddata <= 8'h38;
            14'h1CF0: rddata <= 8'h1E; 14'h1CF1: rddata <= 8'h06; 14'h1CF2: rddata <= 8'h0A; 14'h1CF3: rddata <= 8'hB7;
            14'h1CF4: rddata <= 8'hC8; 14'h1CF5: rddata <= 8'h0A; 14'h1CF6: rddata <= 8'hBE; 14'h1CF7: rddata <= 8'h23;
            14'h1CF8: rddata <= 8'h03; 14'h1CF9: rddata <= 8'hC0; 14'h1CFA: rddata <= 8'h1D; 14'h1CFB: rddata <= 8'h20;
            14'h1CFC: rddata <= 8'hF8; 14'h1CFD: rddata <= 8'hC9; 14'h1CFE: rddata <= 8'h46; 14'h1CFF: rddata <= 8'h6F;
            14'h1D00: rddata <= 8'h75; 14'h1D01: rddata <= 8'h6E; 14'h1D02: rddata <= 8'h64; 14'h1D03: rddata <= 8'h3A;
            14'h1D04: rddata <= 8'h20; 14'h1D05: rddata <= 8'h00; 14'h1D06: rddata <= 8'h53; 14'h1D07: rddata <= 8'h6B;
            14'h1D08: rddata <= 8'h69; 14'h1D09: rddata <= 8'h70; 14'h1D0A: rddata <= 8'h3A; 14'h1D0B: rddata <= 8'h20;
            14'h1D0C: rddata <= 8'h00; 14'h1D0D: rddata <= 8'hD5; 14'h1D0E: rddata <= 8'hF5; 14'h1D0F: rddata <= 8'hCD;
            14'h1D10: rddata <= 8'h9D; 14'h1D11: rddata <= 8'h0E; 14'h1D12: rddata <= 8'h21; 14'h1D13: rddata <= 8'h57;
            14'h1D14: rddata <= 8'h38; 14'h1D15: rddata <= 8'h06; 14'h1D16: rddata <= 8'h06; 14'h1D17: rddata <= 8'h7E;
            14'h1D18: rddata <= 8'h23; 14'h1D19: rddata <= 8'hB7; 14'h1D1A: rddata <= 8'h28; 14'h1D1B: rddata <= 8'h01;
            14'h1D1C: rddata <= 8'hDF; 14'h1D1D: rddata <= 8'h10; 14'h1D1E: rddata <= 8'hF8; 14'h1D1F: rddata <= 8'hCD;
            14'h1D20: rddata <= 8'hEA; 14'h1D21: rddata <= 8'h19; 14'h1D22: rddata <= 8'hF1; 14'h1D23: rddata <= 8'hD1;
            14'h1D24: rddata <= 8'hC9; 14'h1D25: rddata <= 8'hCD; 14'h1D26: rddata <= 8'h7F; 14'h1D27: rddata <= 8'h1B;
            14'h1D28: rddata <= 8'hCD; 14'h1D29: rddata <= 8'hBC; 14'h1D2A: rddata <= 8'h1B; 14'h1D2B: rddata <= 8'h06;
            14'h1D2C: rddata <= 8'h06; 14'h1D2D: rddata <= 8'h21; 14'h1D2E: rddata <= 8'h51; 14'h1D2F: rddata <= 8'h38;
            14'h1D30: rddata <= 8'h7E; 14'h1D31: rddata <= 8'h23; 14'h1D32: rddata <= 8'hCD; 14'h1D33: rddata <= 8'h8A;
            14'h1D34: rddata <= 8'h1B; 14'h1D35: rddata <= 8'h10; 14'h1D36: rddata <= 8'hF9; 14'h1D37: rddata <= 8'hC9;
            14'h1D38: rddata <= 8'hCD; 14'h1D39: rddata <= 8'hBC; 14'h1D3A: rddata <= 8'h1B; 14'h1D3B: rddata <= 8'hEB;
            14'h1D3C: rddata <= 8'h2A; 14'h1D3D: rddata <= 8'hD6; 14'h1D3E: rddata <= 8'h38; 14'h1D3F: rddata <= 8'h1A;
            14'h1D40: rddata <= 8'h13; 14'h1D41: rddata <= 8'hCD; 14'h1D42: rddata <= 8'h8A; 14'h1D43: rddata <= 8'h1B;
            14'h1D44: rddata <= 8'hE7; 14'h1D45: rddata <= 8'h20; 14'h1D46: rddata <= 8'hF8; 14'h1D47: rddata <= 8'hC9;
            14'h1D48: rddata <= 8'h01; 14'h1D49: rddata <= 8'h00; 14'h1D4A: rddata <= 8'h00; 14'h1D4B: rddata <= 8'h0B;
            14'h1D4C: rddata <= 8'h78; 14'h1D4D: rddata <= 8'hB1; 14'h1D4E: rddata <= 8'h20; 14'h1D4F: rddata <= 8'hFB;
            14'h1D50: rddata <= 8'hC9; 14'h1D51: rddata <= 8'hCD; 14'h1D52: rddata <= 8'hCE; 14'h1D53: rddata <= 8'h1B;
            14'h1D54: rddata <= 8'h3E; 14'h1D55: rddata <= 8'hFF; 14'h1D56: rddata <= 8'h32; 14'h1D57: rddata <= 8'h5D;
            14'h1D58: rddata <= 8'h38; 14'h1D59: rddata <= 8'h9F; 14'h1D5A: rddata <= 8'h2F; 14'h1D5B: rddata <= 8'h57;
            14'h1D5C: rddata <= 8'h06; 14'h1D5D: rddata <= 8'h0A; 14'h1D5E: rddata <= 8'hCD; 14'h1D5F: rddata <= 8'h4D;
            14'h1D60: rddata <= 8'h1B; 14'h1D61: rddata <= 8'h5F; 14'h1D62: rddata <= 8'h96; 14'h1D63: rddata <= 8'hA2;
            14'h1D64: rddata <= 8'hC0; 14'h1D65: rddata <= 8'h73; 14'h1D66: rddata <= 8'hCD; 14'h1D67: rddata <= 8'hA9;
            14'h1D68: rddata <= 8'h0B; 14'h1D69: rddata <= 8'h7E; 14'h1D6A: rddata <= 8'hB7; 14'h1D6B: rddata <= 8'h23;
            14'h1D6C: rddata <= 8'h20; 14'h1D6D: rddata <= 8'hEE; 14'h1D6E: rddata <= 8'h10; 14'h1D6F: rddata <= 8'hEE;
            14'h1D70: rddata <= 8'hAF; 14'h1D71: rddata <= 8'hC9; 14'h1D72: rddata <= 8'hF7; 14'h1D73: rddata <= 8'h13;
            14'h1D74: rddata <= 8'hF5; 14'h1D75: rddata <= 8'hFE; 14'h1D76: rddata <= 8'h0A; 14'h1D77: rddata <= 8'h28;
            14'h1D78: rddata <= 8'h1A; 14'h1D79: rddata <= 8'h3A; 14'h1D7A: rddata <= 8'h00; 14'h1D7B: rddata <= 8'h38;
            14'h1D7C: rddata <= 8'hB7; 14'h1D7D: rddata <= 8'h20; 14'h1D7E: rddata <= 8'h14; 14'h1D7F: rddata <= 8'h3A;
            14'h1D80: rddata <= 8'h08; 14'h1D81: rddata <= 8'h38; 14'h1D82: rddata <= 8'hB7; 14'h1D83: rddata <= 8'h28;
            14'h1D84: rddata <= 8'h0E; 14'h1D85: rddata <= 8'h3D; 14'h1D86: rddata <= 8'h32; 14'h1D87: rddata <= 8'h08;
            14'h1D88: rddata <= 8'h38; 14'h1D89: rddata <= 8'h20; 14'h1D8A: rddata <= 8'h08; 14'h1D8B: rddata <= 8'h3E;
            14'h1D8C: rddata <= 8'h17; 14'h1D8D: rddata <= 8'h32; 14'h1D8E: rddata <= 8'h08; 14'h1D8F: rddata <= 8'h38;
            14'h1D90: rddata <= 8'hCD; 14'h1D91: rddata <= 8'h2F; 14'h1D92: rddata <= 8'h1A; 14'h1D93: rddata <= 8'hF1;
            14'h1D94: rddata <= 8'hF5; 14'h1D95: rddata <= 8'hD9; 14'h1D96: rddata <= 8'hFE; 14'h1D97: rddata <= 8'h07;
            14'h1D98: rddata <= 8'hCA; 14'h1D99: rddata <= 8'h14; 14'h1D9A: rddata <= 8'h1E; 14'h1D9B: rddata <= 8'hFE;
            14'h1D9C: rddata <= 8'h0B; 14'h1D9D: rddata <= 8'hCA; 14'h1D9E: rddata <= 8'h45; 14'h1D9F: rddata <= 8'h1E;
            14'h1DA0: rddata <= 8'h5F; 14'h1DA1: rddata <= 8'h2A; 14'h1DA2: rddata <= 8'h01; 14'h1DA3: rddata <= 8'h38;
            14'h1DA4: rddata <= 8'h3A; 14'h1DA5: rddata <= 8'h0D; 14'h1DA6: rddata <= 8'h38; 14'h1DA7: rddata <= 8'h77;
            14'h1DA8: rddata <= 8'h7B; 14'h1DA9: rddata <= 8'hFE; 14'h1DAA: rddata <= 8'h08; 14'h1DAB: rddata <= 8'h28;
            14'h1DAC: rddata <= 8'h30; 14'h1DAD: rddata <= 8'hFE; 14'h1DAE: rddata <= 8'h0D; 14'h1DAF: rddata <= 8'h28;
            14'h1DB0: rddata <= 8'h0D; 14'h1DB1: rddata <= 8'hFE; 14'h1DB2: rddata <= 8'h0A; 14'h1DB3: rddata <= 8'h28;
            14'h1DB4: rddata <= 8'h13; 14'h1DB5: rddata <= 8'h2A; 14'h1DB6: rddata <= 8'h01; 14'h1DB7: rddata <= 8'h38;
            14'h1DB8: rddata <= 8'h77; 14'h1DB9: rddata <= 8'hCD; 14'h1DBA: rddata <= 8'h1F; 14'h1DBB: rddata <= 8'h1E;
            14'h1DBC: rddata <= 8'h18; 14'h1DBD: rddata <= 8'h2C; 14'h1DBE: rddata <= 8'hED; 14'h1DBF: rddata <= 8'h5B;
            14'h1DC0: rddata <= 8'h00; 14'h1DC1: rddata <= 8'h38; 14'h1DC2: rddata <= 8'hAF; 14'h1DC3: rddata <= 8'h57;
            14'h1DC4: rddata <= 8'hED; 14'h1DC5: rddata <= 8'h52; 14'h1DC6: rddata <= 8'h18; 14'h1DC7: rddata <= 8'h1F;
            14'h1DC8: rddata <= 8'h11; 14'h1DC9: rddata <= 8'hC0; 14'h1DCA: rddata <= 8'h33; 14'h1DCB: rddata <= 8'hE7;
            14'h1DCC: rddata <= 8'hD2; 14'h1DCD: rddata <= 8'hD8; 14'h1DCE: rddata <= 8'h1D; 14'h1DCF: rddata <= 8'h11;
            14'h1DD0: rddata <= 8'h28; 14'h1DD1: rddata <= 8'h00; 14'h1DD2: rddata <= 8'h19; 14'h1DD3: rddata <= 8'h22;
            14'h1DD4: rddata <= 8'h01; 14'h1DD5: rddata <= 8'h38; 14'h1DD6: rddata <= 8'h18; 14'h1DD7: rddata <= 8'h12;
            14'h1DD8: rddata <= 8'hCD; 14'h1DD9: rddata <= 8'hFE; 14'h1DDA: rddata <= 8'h1D; 14'h1DDB: rddata <= 8'h18;
            14'h1DDC: rddata <= 8'h0D; 14'h1DDD: rddata <= 8'h3A; 14'h1DDE: rddata <= 8'h00; 14'h1DDF: rddata <= 8'h38;
            14'h1DE0: rddata <= 8'hB7; 14'h1DE1: rddata <= 8'h28; 14'h1DE2: rddata <= 8'h02; 14'h1DE3: rddata <= 8'h2B;
            14'h1DE4: rddata <= 8'h3D; 14'h1DE5: rddata <= 8'h36; 14'h1DE6: rddata <= 8'h20; 14'h1DE7: rddata <= 8'hCD;
            14'h1DE8: rddata <= 8'h3E; 14'h1DE9: rddata <= 8'h1E; 14'h1DEA: rddata <= 8'h2A; 14'h1DEB: rddata <= 8'h01;
            14'h1DEC: rddata <= 8'h38; 14'h1DED: rddata <= 8'h7E; 14'h1DEE: rddata <= 8'h32; 14'h1DEF: rddata <= 8'h0D;
            14'h1DF0: rddata <= 8'h38; 14'h1DF1: rddata <= 8'h36; 14'h1DF2: rddata <= 8'h7F; 14'h1DF3: rddata <= 8'hD9;
            14'h1DF4: rddata <= 8'hF1; 14'h1DF5: rddata <= 8'hC9; 14'h1DF6: rddata <= 8'h2A; 14'h1DF7: rddata <= 8'h01;
            14'h1DF8: rddata <= 8'h38; 14'h1DF9: rddata <= 8'h3A; 14'h1DFA: rddata <= 8'h0D; 14'h1DFB: rddata <= 8'h38;
            14'h1DFC: rddata <= 8'h77; 14'h1DFD: rddata <= 8'hC9; 14'h1DFE: rddata <= 8'h01; 14'h1DFF: rddata <= 8'h98;
            14'h1E00: rddata <= 8'h03; 14'h1E01: rddata <= 8'h11; 14'h1E02: rddata <= 8'h28; 14'h1E03: rddata <= 8'h30;
            14'h1E04: rddata <= 8'h21; 14'h1E05: rddata <= 8'h50; 14'h1E06: rddata <= 8'h30; 14'h1E07: rddata <= 8'hED;
            14'h1E08: rddata <= 8'hB0; 14'h1E09: rddata <= 8'h06; 14'h1E0A: rddata <= 8'h28; 14'h1E0B: rddata <= 8'h21;
            14'h1E0C: rddata <= 8'hC1; 14'h1E0D: rddata <= 8'h33; 14'h1E0E: rddata <= 8'h36; 14'h1E0F: rddata <= 8'h20;
            14'h1E10: rddata <= 8'h23; 14'h1E11: rddata <= 8'h10; 14'h1E12: rddata <= 8'hFB; 14'h1E13: rddata <= 8'hC9;
            14'h1E14: rddata <= 8'h01; 14'h1E15: rddata <= 8'hC8; 14'h1E16: rddata <= 8'h00; 14'h1E17: rddata <= 8'h11;
            14'h1E18: rddata <= 8'h32; 14'h1E19: rddata <= 8'h00; 14'h1E1A: rddata <= 8'hCD; 14'h1E1B: rddata <= 8'h64;
            14'h1E1C: rddata <= 8'h1E; 14'h1E1D: rddata <= 8'h18; 14'h1E1E: rddata <= 8'hD4; 14'h1E1F: rddata <= 8'h2A;
            14'h1E20: rddata <= 8'h01; 14'h1E21: rddata <= 8'h38; 14'h1E22: rddata <= 8'h3A; 14'h1E23: rddata <= 8'h00;
            14'h1E24: rddata <= 8'h38; 14'h1E25: rddata <= 8'h23; 14'h1E26: rddata <= 8'h3C; 14'h1E27: rddata <= 8'hFE;
            14'h1E28: rddata <= 8'h26; 14'h1E29: rddata <= 8'h38; 14'h1E2A: rddata <= 8'h13; 14'h1E2B: rddata <= 8'h23;
            14'h1E2C: rddata <= 8'h23; 14'h1E2D: rddata <= 8'h11; 14'h1E2E: rddata <= 8'hE8; 14'h1E2F: rddata <= 8'h33;
            14'h1E30: rddata <= 8'hE7; 14'h1E31: rddata <= 8'h3E; 14'h1E32: rddata <= 8'h00; 14'h1E33: rddata <= 8'h38;
            14'h1E34: rddata <= 8'h09; 14'h1E35: rddata <= 8'h21; 14'h1E36: rddata <= 8'hC1; 14'h1E37: rddata <= 8'h33;
            14'h1E38: rddata <= 8'hCD; 14'h1E39: rddata <= 8'h3E; 14'h1E3A: rddata <= 8'h1E; 14'h1E3B: rddata <= 8'hC3;
            14'h1E3C: rddata <= 8'hFE; 14'h1E3D: rddata <= 8'h1D; 14'h1E3E: rddata <= 8'h22; 14'h1E3F: rddata <= 8'h01;
            14'h1E40: rddata <= 8'h38; 14'h1E41: rddata <= 8'h32; 14'h1E42: rddata <= 8'h00; 14'h1E43: rddata <= 8'h38;
            14'h1E44: rddata <= 8'hC9; 14'h1E45: rddata <= 8'h06; 14'h1E46: rddata <= 8'h20; 14'h1E47: rddata <= 8'h21;
            14'h1E48: rddata <= 8'h00; 14'h1E49: rddata <= 8'h30; 14'h1E4A: rddata <= 8'hCD; 14'h1E4B: rddata <= 8'h59;
            14'h1E4C: rddata <= 8'h1E; 14'h1E4D: rddata <= 8'h06; 14'h1E4E: rddata <= 8'h06; 14'h1E4F: rddata <= 8'hCD;
            14'h1E50: rddata <= 8'h59; 14'h1E51: rddata <= 8'h1E; 14'h1E52: rddata <= 8'h21; 14'h1E53: rddata <= 8'h29;
            14'h1E54: rddata <= 8'h30; 14'h1E55: rddata <= 8'hAF; 14'h1E56: rddata <= 8'hC3; 14'h1E57: rddata <= 8'hE7;
            14'h1E58: rddata <= 8'h1D; 14'h1E59: rddata <= 8'h11; 14'h1E5A: rddata <= 8'hFF; 14'h1E5B: rddata <= 8'h03;
            14'h1E5C: rddata <= 8'h70; 14'h1E5D: rddata <= 8'h23; 14'h1E5E: rddata <= 8'h1B; 14'h1E5F: rddata <= 8'h7A;
            14'h1E60: rddata <= 8'hB3; 14'h1E61: rddata <= 8'h20; 14'h1E62: rddata <= 8'hF9; 14'h1E63: rddata <= 8'hC9;
            14'h1E64: rddata <= 8'h78; 14'h1E65: rddata <= 8'hB1; 14'h1E66: rddata <= 8'hC8; 14'h1E67: rddata <= 8'hAF;
            14'h1E68: rddata <= 8'hD3; 14'h1E69: rddata <= 8'hFC; 14'h1E6A: rddata <= 8'hCD; 14'h1E6B: rddata <= 8'h76;
            14'h1E6C: rddata <= 8'h1E; 14'h1E6D: rddata <= 8'h3C; 14'h1E6E: rddata <= 8'hD3; 14'h1E6F: rddata <= 8'hFC;
            14'h1E70: rddata <= 8'hCD; 14'h1E71: rddata <= 8'h76; 14'h1E72: rddata <= 8'h1E; 14'h1E73: rddata <= 8'h0B;
            14'h1E74: rddata <= 8'h18; 14'h1E75: rddata <= 8'hEE; 14'h1E76: rddata <= 8'hD5; 14'h1E77: rddata <= 8'hE1;
            14'h1E78: rddata <= 8'h7C; 14'h1E79: rddata <= 8'hB5; 14'h1E7A: rddata <= 8'hC8; 14'h1E7B: rddata <= 8'h2B;
            14'h1E7C: rddata <= 8'h18; 14'h1E7D: rddata <= 8'hFA; 14'h1E7E: rddata <= 8'hF7; 14'h1E7F: rddata <= 8'h12;
            14'h1E80: rddata <= 8'hD9; 14'h1E81: rddata <= 8'h2A; 14'h1E82: rddata <= 8'h0B; 14'h1E83: rddata <= 8'h38;
            14'h1E84: rddata <= 8'h7C; 14'h1E85: rddata <= 8'hB7; 14'h1E86: rddata <= 8'h28; 14'h1E87: rddata <= 8'h1A;
            14'h1E88: rddata <= 8'hEB; 14'h1E89: rddata <= 8'h21; 14'h1E8A: rddata <= 8'h0F; 14'h1E8B: rddata <= 8'h38;
            14'h1E8C: rddata <= 8'h34; 14'h1E8D: rddata <= 8'h7E; 14'h1E8E: rddata <= 8'hFE; 14'h1E8F: rddata <= 8'h0F;
            14'h1E90: rddata <= 8'h38; 14'h1E91: rddata <= 8'h3C; 14'h1E92: rddata <= 8'h36; 14'h1E93: rddata <= 8'h05;
            14'h1E94: rddata <= 8'hEB; 14'h1E95: rddata <= 8'h23; 14'h1E96: rddata <= 8'h7E; 14'h1E97: rddata <= 8'h22;
            14'h1E98: rddata <= 8'h0B; 14'h1E99: rddata <= 8'h38; 14'h1E9A: rddata <= 8'hB7; 14'h1E9B: rddata <= 8'hF2;
            14'h1E9C: rddata <= 8'h36; 14'h1E9D: rddata <= 8'h1F; 14'h1E9E: rddata <= 8'hAF; 14'h1E9F: rddata <= 8'h32;
            14'h1EA0: rddata <= 8'h0C; 14'h1EA1: rddata <= 8'h38; 14'h1EA2: rddata <= 8'h01; 14'h1EA3: rddata <= 8'hFF;
            14'h1EA4: rddata <= 8'h00; 14'h1EA5: rddata <= 8'hED; 14'h1EA6: rddata <= 8'h78; 14'h1EA7: rddata <= 8'h2F;
            14'h1EA8: rddata <= 8'hE6; 14'h1EA9: rddata <= 8'h3F; 14'h1EAA: rddata <= 8'h21; 14'h1EAB: rddata <= 8'h0E;
            14'h1EAC: rddata <= 8'h38; 14'h1EAD: rddata <= 8'h28; 14'h1EAE: rddata <= 8'h16; 14'h1EAF: rddata <= 8'h06;
            14'h1EB0: rddata <= 8'h7F; 14'h1EB1: rddata <= 8'hED; 14'h1EB2: rddata <= 8'h78; 14'h1EB3: rddata <= 8'h2F;
            14'h1EB4: rddata <= 8'hE6; 14'h1EB5: rddata <= 8'h0F; 14'h1EB6: rddata <= 8'h20; 14'h1EB7: rddata <= 8'h1F;
            14'h1EB8: rddata <= 8'h06; 14'h1EB9: rddata <= 8'hBF; 14'h1EBA: rddata <= 8'hED; 14'h1EBB: rddata <= 8'h78;
            14'h1EBC: rddata <= 8'h2F; 14'h1EBD: rddata <= 8'hE6; 14'h1EBE: rddata <= 8'h3F; 14'h1EBF: rddata <= 8'h20;
            14'h1EC0: rddata <= 8'h16; 14'h1EC1: rddata <= 8'hCB; 14'h1EC2: rddata <= 8'h08; 14'h1EC3: rddata <= 8'h38;
            14'h1EC4: rddata <= 8'hF5; 14'h1EC5: rddata <= 8'h23; 14'h1EC6: rddata <= 8'h3E; 14'h1EC7: rddata <= 8'h46;
            14'h1EC8: rddata <= 8'hBE; 14'h1EC9: rddata <= 8'h38; 14'h1ECA: rddata <= 8'h03; 14'h1ECB: rddata <= 8'h28;
            14'h1ECC: rddata <= 8'h04; 14'h1ECD: rddata <= 8'h34; 14'h1ECE: rddata <= 8'hAF; 14'h1ECF: rddata <= 8'hD9;
            14'h1ED0: rddata <= 8'hC9; 14'h1ED1: rddata <= 8'h34; 14'h1ED2: rddata <= 8'h2B; 14'h1ED3: rddata <= 8'h36;
            14'h1ED4: rddata <= 8'h00; 14'h1ED5: rddata <= 8'h18; 14'h1ED6: rddata <= 8'hF7; 14'h1ED7: rddata <= 8'h11;
            14'h1ED8: rddata <= 8'h00; 14'h1ED9: rddata <= 8'h00; 14'h1EDA: rddata <= 8'h1C; 14'h1EDB: rddata <= 8'h1F;
            14'h1EDC: rddata <= 8'h30; 14'h1EDD: rddata <= 8'hFC; 14'h1EDE: rddata <= 8'h7B; 14'h1EDF: rddata <= 8'hCB;
            14'h1EE0: rddata <= 8'h18; 14'h1EE1: rddata <= 8'h30; 14'h1EE2: rddata <= 8'h04; 14'h1EE3: rddata <= 8'hC6;
            14'h1EE4: rddata <= 8'h06; 14'h1EE5: rddata <= 8'h18; 14'h1EE6: rddata <= 8'hF8; 14'h1EE7: rddata <= 8'h5F;
            14'h1EE8: rddata <= 8'hBE; 14'h1EE9: rddata <= 8'h77; 14'h1EEA: rddata <= 8'h23; 14'h1EEB: rddata <= 8'h20;
            14'h1EEC: rddata <= 8'h0F; 14'h1EED: rddata <= 8'h3E; 14'h1EEE: rddata <= 8'h04; 14'h1EEF: rddata <= 8'hBE;
            14'h1EF0: rddata <= 8'h38; 14'h1EF1: rddata <= 8'h05; 14'h1EF2: rddata <= 8'h28; 14'h1EF3: rddata <= 8'h0C;
            14'h1EF4: rddata <= 8'h34; 14'h1EF5: rddata <= 8'h18; 14'h1EF6: rddata <= 8'h02; 14'h1EF7: rddata <= 8'h36;
            14'h1EF8: rddata <= 8'h06; 14'h1EF9: rddata <= 8'hAF; 14'h1EFA: rddata <= 8'hD9; 14'h1EFB: rddata <= 8'hC9;
            14'h1EFC: rddata <= 8'h36; 14'h1EFD: rddata <= 8'h00; 14'h1EFE: rddata <= 8'h18; 14'h1EFF: rddata <= 8'hF9;
            14'h1F00: rddata <= 8'h34; 14'h1F01: rddata <= 8'h06; 14'h1F02: rddata <= 8'h7F; 14'h1F03: rddata <= 8'hED;
            14'h1F04: rddata <= 8'h78; 14'h1F05: rddata <= 8'hCB; 14'h1F06: rddata <= 8'h6F; 14'h1F07: rddata <= 8'hDD;
            14'h1F08: rddata <= 8'h21; 14'h1F09: rddata <= 8'h93; 14'h1F0A: rddata <= 8'h1F; 14'h1F0B: rddata <= 8'h28;
            14'h1F0C: rddata <= 8'h0C; 14'h1F0D: rddata <= 8'hCB; 14'h1F0E: rddata <= 8'h67; 14'h1F0F: rddata <= 8'hDD;
            14'h1F10: rddata <= 8'h21; 14'h1F11: rddata <= 8'h65; 14'h1F12: rddata <= 8'h1F; 14'h1F13: rddata <= 8'h28;
            14'h1F14: rddata <= 8'h04; 14'h1F15: rddata <= 8'hDD; 14'h1F16: rddata <= 8'h21; 14'h1F17: rddata <= 8'h37;
            14'h1F18: rddata <= 8'h1F; 14'h1F19: rddata <= 8'hDD; 14'h1F1A: rddata <= 8'h19; 14'h1F1B: rddata <= 8'hDD;
            14'h1F1C: rddata <= 8'h7E; 14'h1F1D: rddata <= 8'h00; 14'h1F1E: rddata <= 8'hB7; 14'h1F1F: rddata <= 8'hF2;
            14'h1F20: rddata <= 8'h36; 14'h1F21: rddata <= 8'h1F; 14'h1F22: rddata <= 8'hD6; 14'h1F23: rddata <= 8'h7F;
            14'h1F24: rddata <= 8'h4F; 14'h1F25: rddata <= 8'h21; 14'h1F26: rddata <= 8'h44; 14'h1F27: rddata <= 8'h02;
            14'h1F28: rddata <= 8'h23; 14'h1F29: rddata <= 8'h7E; 14'h1F2A: rddata <= 8'hB7; 14'h1F2B: rddata <= 8'hF2;
            14'h1F2C: rddata <= 8'h28; 14'h1F2D: rddata <= 8'h1F; 14'h1F2E: rddata <= 8'h0D; 14'h1F2F: rddata <= 8'h20;
            14'h1F30: rddata <= 8'hF7; 14'h1F31: rddata <= 8'h22; 14'h1F32: rddata <= 8'h0B; 14'h1F33: rddata <= 8'h38;
            14'h1F34: rddata <= 8'hE6; 14'h1F35: rddata <= 8'h7F; 14'h1F36: rddata <= 8'hD9; 14'h1F37: rddata <= 8'hC9;
            14'h1F38: rddata <= 8'h3D; 14'h1F39: rddata <= 8'h08; 14'h1F3A: rddata <= 8'h3A; 14'h1F3B: rddata <= 8'h0D;
            14'h1F3C: rddata <= 8'h3B; 14'h1F3D: rddata <= 8'h2E; 14'h1F3E: rddata <= 8'h2D; 14'h1F3F: rddata <= 8'h2F;
            14'h1F40: rddata <= 8'h30; 14'h1F41: rddata <= 8'h70; 14'h1F42: rddata <= 8'h6C; 14'h1F43: rddata <= 8'h2C;
            14'h1F44: rddata <= 8'h39; 14'h1F45: rddata <= 8'h6F; 14'h1F46: rddata <= 8'h6B; 14'h1F47: rddata <= 8'h6D;
            14'h1F48: rddata <= 8'h6E; 14'h1F49: rddata <= 8'h6A; 14'h1F4A: rddata <= 8'h38; 14'h1F4B: rddata <= 8'h69;
            14'h1F4C: rddata <= 8'h37; 14'h1F4D: rddata <= 8'h75; 14'h1F4E: rddata <= 8'h68; 14'h1F4F: rddata <= 8'h62;
            14'h1F50: rddata <= 8'h36; 14'h1F51: rddata <= 8'h79; 14'h1F52: rddata <= 8'h67; 14'h1F53: rddata <= 8'h76;
            14'h1F54: rddata <= 8'h63; 14'h1F55: rddata <= 8'h66; 14'h1F56: rddata <= 8'h35; 14'h1F57: rddata <= 8'h74;
            14'h1F58: rddata <= 8'h34; 14'h1F59: rddata <= 8'h72; 14'h1F5A: rddata <= 8'h64; 14'h1F5B: rddata <= 8'h78;
            14'h1F5C: rddata <= 8'h33; 14'h1F5D: rddata <= 8'h65; 14'h1F5E: rddata <= 8'h73; 14'h1F5F: rddata <= 8'h7A;
            14'h1F60: rddata <= 8'h20; 14'h1F61: rddata <= 8'h61; 14'h1F62: rddata <= 8'h32; 14'h1F63: rddata <= 8'h77;
            14'h1F64: rddata <= 8'h31; 14'h1F65: rddata <= 8'h71; 14'h1F66: rddata <= 8'h2B; 14'h1F67: rddata <= 8'h5C;
            14'h1F68: rddata <= 8'h2A; 14'h1F69: rddata <= 8'h0D; 14'h1F6A: rddata <= 8'h40; 14'h1F6B: rddata <= 8'h3E;
            14'h1F6C: rddata <= 8'h5F; 14'h1F6D: rddata <= 8'h5E; 14'h1F6E: rddata <= 8'h3F; 14'h1F6F: rddata <= 8'h50;
            14'h1F70: rddata <= 8'h4C; 14'h1F71: rddata <= 8'h3C; 14'h1F72: rddata <= 8'h29; 14'h1F73: rddata <= 8'h4F;
            14'h1F74: rddata <= 8'h4B; 14'h1F75: rddata <= 8'h4D; 14'h1F76: rddata <= 8'h4E; 14'h1F77: rddata <= 8'h4A;
            14'h1F78: rddata <= 8'h28; 14'h1F79: rddata <= 8'h49; 14'h1F7A: rddata <= 8'h27; 14'h1F7B: rddata <= 8'h55;
            14'h1F7C: rddata <= 8'h48; 14'h1F7D: rddata <= 8'h42; 14'h1F7E: rddata <= 8'h26; 14'h1F7F: rddata <= 8'h59;
            14'h1F80: rddata <= 8'h47; 14'h1F81: rddata <= 8'h56; 14'h1F82: rddata <= 8'h43; 14'h1F83: rddata <= 8'h46;
            14'h1F84: rddata <= 8'h25; 14'h1F85: rddata <= 8'h54; 14'h1F86: rddata <= 8'h24; 14'h1F87: rddata <= 8'h52;
            14'h1F88: rddata <= 8'h44; 14'h1F89: rddata <= 8'h58; 14'h1F8A: rddata <= 8'h23; 14'h1F8B: rddata <= 8'h45;
            14'h1F8C: rddata <= 8'h53; 14'h1F8D: rddata <= 8'h5A; 14'h1F8E: rddata <= 8'h20; 14'h1F8F: rddata <= 8'h41;
            14'h1F90: rddata <= 8'h22; 14'h1F91: rddata <= 8'h57; 14'h1F92: rddata <= 8'h21; 14'h1F93: rddata <= 8'h51;
            14'h1F94: rddata <= 8'h82; 14'h1F95: rddata <= 8'h1C; 14'h1F96: rddata <= 8'hC1; 14'h1F97: rddata <= 8'h0D;
            14'h1F98: rddata <= 8'h94; 14'h1F99: rddata <= 8'hC4; 14'h1F9A: rddata <= 8'h81; 14'h1F9B: rddata <= 8'h1E;
            14'h1F9C: rddata <= 8'h30; 14'h1F9D: rddata <= 8'h10; 14'h1F9E: rddata <= 8'hCA; 14'h1F9F: rddata <= 8'hC3;
            14'h1FA0: rddata <= 8'h92; 14'h1FA1: rddata <= 8'h0F; 14'h1FA2: rddata <= 8'h9D; 14'h1FA3: rddata <= 8'h0D;
            14'h1FA4: rddata <= 8'hC8; 14'h1FA5: rddata <= 8'h9C; 14'h1FA6: rddata <= 8'h8D; 14'h1FA7: rddata <= 8'h09;
            14'h1FA8: rddata <= 8'h8C; 14'h1FA9: rddata <= 8'h15; 14'h1FAA: rddata <= 8'h08; 14'h1FAB: rddata <= 8'hC9;
            14'h1FAC: rddata <= 8'h90; 14'h1FAD: rddata <= 8'h19; 14'h1FAE: rddata <= 8'h07; 14'h1FAF: rddata <= 8'hC7;
            14'h1FB0: rddata <= 8'h03; 14'h1FB1: rddata <= 8'h83; 14'h1FB2: rddata <= 8'h88; 14'h1FB3: rddata <= 8'h84;
            14'h1FB4: rddata <= 8'hA5; 14'h1FB5: rddata <= 8'h12; 14'h1FB6: rddata <= 8'h86; 14'h1FB7: rddata <= 8'h18;
            14'h1FB8: rddata <= 8'h8A; 14'h1FB9: rddata <= 8'h85; 14'h1FBA: rddata <= 8'h13; 14'h1FBB: rddata <= 8'h9A;
            14'h1FBC: rddata <= 8'hC6; 14'h1FBD: rddata <= 8'h9B; 14'h1FBE: rddata <= 8'h97; 14'h1FBF: rddata <= 8'h8E;
            14'h1FC0: rddata <= 8'h89; 14'h1FC1: rddata <= 8'h11; 14'h1FC2: rddata <= 8'hE5; 14'h1FC3: rddata <= 8'h21;
            14'h1FC4: rddata <= 8'h04; 14'h1FC5: rddata <= 8'h00; 14'h1FC6: rddata <= 8'h39; 14'h1FC7: rddata <= 8'h22;
            14'h1FC8: rddata <= 8'hF9; 14'h1FC9: rddata <= 8'h38; 14'h1FCA: rddata <= 8'hE1; 14'h1FCB: rddata <= 8'hC3;
            14'h1FCC: rddata <= 8'h25; 14'h1FCD: rddata <= 8'h1A; 14'h1FCE: rddata <= 8'h2A; 14'h1FCF: rddata <= 8'hF9;
            14'h1FD0: rddata <= 8'h38; 14'h1FD1: rddata <= 8'hF9; 14'h1FD2: rddata <= 8'h2A; 14'h1FD3: rddata <= 8'hCE;
            14'h1FD4: rddata <= 8'h38; 14'h1FD5: rddata <= 8'hCD; 14'h1FD6: rddata <= 8'h20; 14'h1FD7: rddata <= 8'h0C;
            14'h1FD8: rddata <= 8'h2B; 14'h1FD9: rddata <= 8'h2B; 14'h1FDA: rddata <= 8'h22; 14'h1FDB: rddata <= 8'hF9;
            14'h1FDC: rddata <= 8'h38; 14'h1FDD: rddata <= 8'h21; 14'h1FDE: rddata <= 8'hB1; 14'h1FDF: rddata <= 8'h38;
            14'h1FE0: rddata <= 8'hC9; 14'h1FE1: rddata <= 8'h3E; 14'h1FE2: rddata <= 8'hFF; 14'h1FE3: rddata <= 8'hD3;
            14'h1FE4: rddata <= 8'hFE; 14'h1FE5: rddata <= 8'hC3; 14'h1FE6: rddata <= 8'h41; 14'h1FE7: rddata <= 8'h00;
            14'h1FE8: rddata <= 8'h3E; 14'h1FE9: rddata <= 8'hAA; 14'h1FEA: rddata <= 8'hD3; 14'h1FEB: rddata <= 8'hFF;
            14'h1FEC: rddata <= 8'h32; 14'h1FED: rddata <= 8'h09; 14'h1FEE: rddata <= 8'h38; 14'h1FEF: rddata <= 8'hC3;
            14'h1FF0: rddata <= 8'h10; 14'h1FF1: rddata <= 8'h20; 14'h1FF2: rddata <= 8'h21; 14'h1FF3: rddata <= 8'h5F;
            14'h1FF4: rddata <= 8'h01; 14'h1FF5: rddata <= 8'hC3; 14'h1FF6: rddata <= 8'h9D; 14'h1FF7: rddata <= 8'h0E;
            14'h1FF8: rddata <= 8'hF5; 14'h1FF9: rddata <= 8'hF5; 14'h1FFA: rddata <= 8'hF5; 14'h1FFB: rddata <= 8'hF5;
            14'h1FFC: rddata <= 8'hF5; 14'h1FFD: rddata <= 8'hF5; 14'h1FFE: rddata <= 8'hF5; 14'h1FFF: rddata <= 8'hF5;
            14'h2000: rddata <= 8'hC3; 14'h2001: rddata <= 8'h09; 14'h2002: rddata <= 8'h20; 14'h2003: rddata <= 8'hC3;
            14'h2004: rddata <= 8'h7E; 14'h2005: rddata <= 8'h20; 14'h2006: rddata <= 8'hC3; 14'h2007: rddata <= 8'hD3;
            14'h2008: rddata <= 8'h20; 14'h2009: rddata <= 8'h31; 14'h200A: rddata <= 8'hA0; 14'h200B: rddata <= 8'h38;
            14'h200C: rddata <= 8'h3E; 14'h200D: rddata <= 8'hC0; 14'h200E: rddata <= 8'hD3; 14'h200F: rddata <= 8'hF0;
            14'h2010: rddata <= 8'h3E; 14'h2011: rddata <= 8'h21; 14'h2012: rddata <= 8'hD3; 14'h2013: rddata <= 8'hF1;
            14'h2014: rddata <= 8'h3E; 14'h2015: rddata <= 8'h22; 14'h2016: rddata <= 8'hD3; 14'h2017: rddata <= 8'hF2;
            14'h2018: rddata <= 8'h3E; 14'h2019: rddata <= 8'h13; 14'h201A: rddata <= 8'hD3; 14'h201B: rddata <= 8'hF3;
            14'h201C: rddata <= 8'h3E; 14'h201D: rddata <= 8'h01; 14'h201E: rddata <= 8'hD3; 14'h201F: rddata <= 8'hE0;
            14'h2020: rddata <= 8'h21; 14'h2021: rddata <= 8'h3E; 14'h2022: rddata <= 8'h20; 14'h2023: rddata <= 8'h0E;
            14'h2024: rddata <= 8'hEA; 14'h2025: rddata <= 8'h06; 14'h2026: rddata <= 8'h00; 14'h2027: rddata <= 8'h16;
            14'h2028: rddata <= 8'h20; 14'h2029: rddata <= 8'hED; 14'h202A: rddata <= 8'h41; 14'h202B: rddata <= 8'h7E;
            14'h202C: rddata <= 8'hD3; 14'h202D: rddata <= 8'hEB; 14'h202E: rddata <= 8'h23; 14'h202F: rddata <= 8'h04;
            14'h2030: rddata <= 8'h15; 14'h2031: rddata <= 8'h20; 14'h2032: rddata <= 8'hF6; 14'h2033: rddata <= 8'hCD;
            14'h2034: rddata <= 8'h5E; 14'h2035: rddata <= 8'h20; 14'h2036: rddata <= 8'h3E; 14'h2037: rddata <= 8'h01;
            14'h2038: rddata <= 8'hCD; 14'h2039: rddata <= 8'hEF; 14'h203A: rddata <= 8'h25; 14'h203B: rddata <= 8'hC3;
            14'h203C: rddata <= 8'hE1; 14'h203D: rddata <= 8'h1F; 14'h203E: rddata <= 8'h11; 14'h203F: rddata <= 8'h01;
            14'h2040: rddata <= 8'h11; 14'h2041: rddata <= 8'h0F; 14'h2042: rddata <= 8'hF1; 14'h2043: rddata <= 8'h01;
            14'h2044: rddata <= 8'hF1; 14'h2045: rddata <= 8'h0F; 14'h2046: rddata <= 8'h2E; 14'h2047: rddata <= 8'h02;
            14'h2048: rddata <= 8'h1F; 14'h2049: rddata <= 8'h0F; 14'h204A: rddata <= 8'hCC; 14'h204B: rddata <= 8'h03;
            14'h204C: rddata <= 8'hFF; 14'h204D: rddata <= 8'h0F; 14'h204E: rddata <= 8'hCC; 14'h204F: rddata <= 8'h0C;
            14'h2050: rddata <= 8'hBB; 14'h2051: rddata <= 8'h03; 14'h2052: rddata <= 8'h2C; 14'h2053: rddata <= 8'h0C;
            14'h2054: rddata <= 8'h19; 14'h2055: rddata <= 8'h04; 14'h2056: rddata <= 8'hF7; 14'h2057: rddata <= 8'h0F;
            14'h2058: rddata <= 8'hD4; 14'h2059: rddata <= 8'h02; 14'h205A: rddata <= 8'h22; 14'h205B: rddata <= 8'h0B;
            14'h205C: rddata <= 8'h33; 14'h205D: rddata <= 8'h03; 14'h205E: rddata <= 8'hDB; 14'h205F: rddata <= 8'hF1;
            14'h2060: rddata <= 8'hF5; 14'h2061: rddata <= 8'hDB; 14'h2062: rddata <= 8'hF2; 14'h2063: rddata <= 8'hF5;
            14'h2064: rddata <= 8'h3E; 14'h2065: rddata <= 8'h15; 14'h2066: rddata <= 8'hD3; 14'h2067: rddata <= 8'hF1;
            14'h2068: rddata <= 8'h3E; 14'h2069: rddata <= 8'h00; 14'h206A: rddata <= 8'hD3; 14'h206B: rddata <= 8'hF2;
            14'h206C: rddata <= 8'h11; 14'h206D: rddata <= 8'h00; 14'h206E: rddata <= 8'h40; 14'h206F: rddata <= 8'h21;
            14'h2070: rddata <= 8'h00; 14'h2071: rddata <= 8'hB0; 14'h2072: rddata <= 8'h01; 14'h2073: rddata <= 8'h00;
            14'h2074: rddata <= 8'h08; 14'h2075: rddata <= 8'hED; 14'h2076: rddata <= 8'hB0; 14'h2077: rddata <= 8'hF1;
            14'h2078: rddata <= 8'hD3; 14'h2079: rddata <= 8'hF2; 14'h207A: rddata <= 8'hF1; 14'h207B: rddata <= 8'hD3;
            14'h207C: rddata <= 8'hF1; 14'h207D: rddata <= 8'hC9; 14'h207E: rddata <= 8'h21; 14'h207F: rddata <= 8'hFF;
            14'h2080: rddata <= 8'hBE; 14'h2081: rddata <= 8'h22; 14'h2082: rddata <= 8'hAD; 14'h2083: rddata <= 8'h38;
            14'h2084: rddata <= 8'h11; 14'h2085: rddata <= 8'hCE; 14'h2086: rddata <= 8'hFF; 14'h2087: rddata <= 8'h19;
            14'h2088: rddata <= 8'h22; 14'h2089: rddata <= 8'h4B; 14'h208A: rddata <= 8'h38; 14'h208B: rddata <= 8'h21;
            14'h208C: rddata <= 8'h00; 14'h208D: rddata <= 8'h39; 14'h208E: rddata <= 8'h36; 14'h208F: rddata <= 8'h00;
            14'h2090: rddata <= 8'h23; 14'h2091: rddata <= 8'h22; 14'h2092: rddata <= 8'h4F; 14'h2093: rddata <= 8'h38;
            14'h2094: rddata <= 8'hCD; 14'h2095: rddata <= 8'hBE; 14'h2096: rddata <= 8'h0B; 14'h2097: rddata <= 8'h21;
            14'h2098: rddata <= 8'hF1; 14'h2099: rddata <= 8'h20; 14'h209A: rddata <= 8'h22; 14'h209B: rddata <= 8'h06;
            14'h209C: rddata <= 8'h38; 14'h209D: rddata <= 8'hCD; 14'h209E: rddata <= 8'hF2; 14'h209F: rddata <= 8'h1F;
            14'h20A0: rddata <= 8'h21; 14'h20A1: rddata <= 8'hBF; 14'h20A2: rddata <= 8'h20; 14'h20A3: rddata <= 8'hCD;
            14'h20A4: rddata <= 8'h9D; 14'h20A5: rddata <= 8'h0E; 14'h20A6: rddata <= 8'h3E; 14'h20A7: rddata <= 8'h02;
            14'h20A8: rddata <= 8'hCD; 14'h20A9: rddata <= 8'hEF; 14'h20AA: rddata <= 8'h25; 14'h20AB: rddata <= 8'hCD;
            14'h20AC: rddata <= 8'h02; 14'h20AD: rddata <= 8'h26; 14'h20AE: rddata <= 8'hB7; 14'h20AF: rddata <= 8'h28;
            14'h20B0: rddata <= 8'h05; 14'h20B1: rddata <= 8'hCD; 14'h20B2: rddata <= 8'h72; 14'h20B3: rddata <= 8'h1D;
            14'h20B4: rddata <= 8'h18; 14'h20B5: rddata <= 8'hF5; 14'h20B6: rddata <= 8'hCD; 14'h20B7: rddata <= 8'hEA;
            14'h20B8: rddata <= 8'h19; 14'h20B9: rddata <= 8'hCD; 14'h20BA: rddata <= 8'hEA; 14'h20BB: rddata <= 8'h19;
            14'h20BC: rddata <= 8'hC3; 14'h20BD: rddata <= 8'h53; 14'h20BE: rddata <= 8'h01; 14'h20BF: rddata <= 8'h0D;
            14'h20C0: rddata <= 8'h0A; 14'h20C1: rddata <= 8'h41; 14'h20C2: rddata <= 8'h71; 14'h20C3: rddata <= 8'h75;
            14'h20C4: rddata <= 8'h61; 14'h20C5: rddata <= 8'h72; 14'h20C6: rddata <= 8'h69; 14'h20C7: rddata <= 8'h75;
            14'h20C8: rddata <= 8'h73; 14'h20C9: rddata <= 8'h2B; 14'h20CA: rddata <= 8'h20; 14'h20CB: rddata <= 8'h53;
            14'h20CC: rddata <= 8'h79; 14'h20CD: rddata <= 8'h73; 14'h20CE: rddata <= 8'h74; 14'h20CF: rddata <= 8'h65;
            14'h20D0: rddata <= 8'h6D; 14'h20D1: rddata <= 8'h20; 14'h20D2: rddata <= 8'h00; 14'h20D3: rddata <= 8'hFE;
            14'h20D4: rddata <= 8'h00; 14'h20D5: rddata <= 8'hC2; 14'h20D6: rddata <= 8'hDB; 14'h20D7: rddata <= 8'h20;
            14'h20D8: rddata <= 8'hC3; 14'h20D9: rddata <= 8'h10; 14'h20DA: rddata <= 8'hE0; 14'h20DB: rddata <= 8'h3E;
            14'h20DC: rddata <= 8'h23; 14'h20DD: rddata <= 8'hD3; 14'h20DE: rddata <= 8'hF2; 14'h20DF: rddata <= 8'h11;
            14'h20E0: rddata <= 8'h00; 14'h20E1: rddata <= 8'h80; 14'h20E2: rddata <= 8'h21; 14'h20E3: rddata <= 8'h00;
            14'h20E4: rddata <= 8'hC0; 14'h20E5: rddata <= 8'h01; 14'h20E6: rddata <= 8'h00; 14'h20E7: rddata <= 8'h40;
            14'h20E8: rddata <= 8'hED; 14'h20E9: rddata <= 8'hB0; 14'h20EA: rddata <= 8'h3E; 14'h20EB: rddata <= 8'h23;
            14'h20EC: rddata <= 8'hD3; 14'h20ED: rddata <= 8'hF3; 14'h20EE: rddata <= 8'hC3; 14'h20EF: rddata <= 8'hF9;
            14'h20F0: rddata <= 8'h28; 14'h20F1: rddata <= 8'hE3; 14'h20F2: rddata <= 8'hF5; 14'h20F3: rddata <= 8'h7E;
            14'h20F4: rddata <= 8'h23; 14'h20F5: rddata <= 8'hE5; 14'h20F6: rddata <= 8'h21; 14'h20F7: rddata <= 8'h13;
            14'h20F8: rddata <= 8'h21; 14'h20F9: rddata <= 8'hC5; 14'h20FA: rddata <= 8'h01; 14'h20FB: rddata <= 8'h06;
            14'h20FC: rddata <= 8'h00; 14'h20FD: rddata <= 8'hED; 14'h20FE: rddata <= 8'hB1; 14'h20FF: rddata <= 8'h79;
            14'h2100: rddata <= 8'hC1; 14'h2101: rddata <= 8'h87; 14'h2102: rddata <= 8'h21; 14'h2103: rddata <= 8'h18;
            14'h2104: rddata <= 8'h21; 14'h2105: rddata <= 8'h85; 14'h2106: rddata <= 8'h6F; 14'h2107: rddata <= 8'hAF;
            14'h2108: rddata <= 8'h8C; 14'h2109: rddata <= 8'h67; 14'h210A: rddata <= 8'h7E; 14'h210B: rddata <= 8'h23;
            14'h210C: rddata <= 8'h66; 14'h210D: rddata <= 8'h6F; 14'h210E: rddata <= 8'hE9; 14'h210F: rddata <= 8'hE1;
            14'h2110: rddata <= 8'hF1; 14'h2111: rddata <= 8'hE3; 14'h2112: rddata <= 8'hC9; 14'h2113: rddata <= 8'h18;
            14'h2114: rddata <= 8'h17; 14'h2115: rddata <= 8'h16; 14'h2116: rddata <= 8'h0A; 14'h2117: rddata <= 8'h1B;
            14'h2118: rddata <= 8'h0F; 14'h2119: rddata <= 8'h21; 14'h211A: rddata <= 8'h7F; 14'h211B: rddata <= 8'h21;
            14'h211C: rddata <= 8'h93; 14'h211D: rddata <= 8'h21; 14'h211E: rddata <= 8'hA6; 14'h211F: rddata <= 8'h21;
            14'h2120: rddata <= 8'hB8; 14'h2121: rddata <= 8'h21; 14'h2122: rddata <= 8'hD4; 14'h2123: rddata <= 8'h21;
            14'h2124: rddata <= 8'hC5; 14'h2125: rddata <= 8'h44; 14'h2126: rddata <= 8'h49; 14'h2127: rddata <= 8'h54;
            14'h2128: rddata <= 8'hC3; 14'h2129: rddata <= 8'h4C; 14'h212A: rddata <= 8'h53; 14'h212B: rddata <= 8'hCC;
            14'h212C: rddata <= 8'h4F; 14'h212D: rddata <= 8'h43; 14'h212E: rddata <= 8'h41; 14'h212F: rddata <= 8'h54;
            14'h2130: rddata <= 8'h45; 14'h2131: rddata <= 8'hCF; 14'h2132: rddata <= 8'h55; 14'h2133: rddata <= 8'h54;
            14'h2134: rddata <= 8'hD0; 14'h2135: rddata <= 8'h53; 14'h2136: rddata <= 8'h47; 14'h2137: rddata <= 8'hC4;
            14'h2138: rddata <= 8'h45; 14'h2139: rddata <= 8'h42; 14'h213A: rddata <= 8'h55; 14'h213B: rddata <= 8'h47;
            14'h213C: rddata <= 8'hC3; 14'h213D: rddata <= 8'h41; 14'h213E: rddata <= 8'h4C; 14'h213F: rddata <= 8'h4C;
            14'h2140: rddata <= 8'hCC; 14'h2141: rddata <= 8'h4F; 14'h2142: rddata <= 8'h41; 14'h2143: rddata <= 8'h44;
            14'h2144: rddata <= 8'hD3; 14'h2145: rddata <= 8'h41; 14'h2146: rddata <= 8'h56; 14'h2147: rddata <= 8'h45;
            14'h2148: rddata <= 8'hC4; 14'h2149: rddata <= 8'h49; 14'h214A: rddata <= 8'h52; 14'h214B: rddata <= 8'hCD;
            14'h214C: rddata <= 8'h4B; 14'h214D: rddata <= 8'h44; 14'h214E: rddata <= 8'h49; 14'h214F: rddata <= 8'h52;
            14'h2150: rddata <= 8'hC4; 14'h2151: rddata <= 8'h45; 14'h2152: rddata <= 8'h4C; 14'h2153: rddata <= 8'hC3;
            14'h2154: rddata <= 8'h44; 14'h2155: rddata <= 8'hC9; 14'h2156: rddata <= 8'h4E; 14'h2157: rddata <= 8'hCA;
            14'h2158: rddata <= 8'h4F; 14'h2159: rddata <= 8'h59; 14'h215A: rddata <= 8'hC8; 14'h215B: rddata <= 8'h45;
            14'h215C: rddata <= 8'h58; 14'h215D: rddata <= 8'h24; 14'h215E: rddata <= 8'h80; 14'h215F: rddata <= 8'hEF;
            14'h2160: rddata <= 8'h21; 14'h2161: rddata <= 8'hF0; 14'h2162: rddata <= 8'h21; 14'h2163: rddata <= 8'h04;
            14'h2164: rddata <= 8'h22; 14'h2165: rddata <= 8'hF4; 14'h2166: rddata <= 8'h21; 14'h2167: rddata <= 8'h43;
            14'h2168: rddata <= 8'h22; 14'h2169: rddata <= 8'hEF; 14'h216A: rddata <= 8'h21; 14'h216B: rddata <= 8'hFC;
            14'h216C: rddata <= 8'h22; 14'h216D: rddata <= 8'h04; 14'h216E: rddata <= 8'h23; 14'h216F: rddata <= 8'h53;
            14'h2170: rddata <= 8'h23; 14'h2171: rddata <= 8'hDE; 14'h2172: rddata <= 8'h23; 14'h2173: rddata <= 8'hCD;
            14'h2174: rddata <= 8'h23; 14'h2175: rddata <= 8'h8E; 14'h2176: rddata <= 8'h23; 14'h2177: rddata <= 8'h9F;
            14'h2178: rddata <= 8'h23; 14'h2179: rddata <= 8'h6C; 14'h217A: rddata <= 8'h22; 14'h217B: rddata <= 8'h80;
            14'h217C: rddata <= 8'h22; 14'h217D: rddata <= 8'hC2; 14'h217E: rddata <= 8'h22; 14'h217F: rddata <= 8'hC1;
            14'h2180: rddata <= 8'hF1; 14'h2181: rddata <= 8'hE1; 14'h2182: rddata <= 8'hC5; 14'h2183: rddata <= 8'hFE;
            14'h2184: rddata <= 8'h2F; 14'h2185: rddata <= 8'hD8; 14'h2186: rddata <= 8'hFE; 14'h2187: rddata <= 8'h32;
            14'h2188: rddata <= 8'hD0; 14'h2189: rddata <= 8'hD6; 14'h218A: rddata <= 8'h2F; 14'h218B: rddata <= 8'h87;
            14'h218C: rddata <= 8'hE5; 14'h218D: rddata <= 8'h21; 14'h218E: rddata <= 8'h79; 14'h218F: rddata <= 8'h21;
            14'h2190: rddata <= 8'hC3; 14'h2191: rddata <= 8'h05; 14'h2192: rddata <= 8'h21; 14'h2193: rddata <= 8'h78;
            14'h2194: rddata <= 8'hFE; 14'h2195: rddata <= 8'hCB; 14'h2196: rddata <= 8'hC2; 14'h2197: rddata <= 8'h0F;
            14'h2198: rddata <= 8'h21; 14'h2199: rddata <= 8'hC1; 14'h219A: rddata <= 8'hF1; 14'h219B: rddata <= 8'hE1;
            14'h219C: rddata <= 8'hC5; 14'h219D: rddata <= 8'hEB; 14'h219E: rddata <= 8'h11; 14'h219F: rddata <= 8'h23;
            14'h21A0: rddata <= 8'h21; 14'h21A1: rddata <= 8'h06; 14'h21A2: rddata <= 8'hD3; 14'h21A3: rddata <= 8'hC3;
            14'h21A4: rddata <= 8'hF9; 14'h21A5: rddata <= 8'h04; 14'h21A6: rddata <= 8'hD1; 14'h21A7: rddata <= 8'hF1;
            14'h21A8: rddata <= 8'hE1; 14'h21A9: rddata <= 8'hFE; 14'h21AA: rddata <= 8'hD4; 14'h21AB: rddata <= 8'h30;
            14'h21AC: rddata <= 8'h02; 14'h21AD: rddata <= 8'hD5; 14'h21AE: rddata <= 8'hC9; 14'h21AF: rddata <= 8'hD6;
            14'h21B0: rddata <= 8'hD3; 14'h21B1: rddata <= 8'h4F; 14'h21B2: rddata <= 8'h11; 14'h21B3: rddata <= 8'h24;
            14'h21B4: rddata <= 8'h21; 14'h21B5: rddata <= 8'hC3; 14'h21B6: rddata <= 8'hA8; 14'h21B7: rddata <= 8'h05;
            14'h21B8: rddata <= 8'hC1; 14'h21B9: rddata <= 8'hF1; 14'h21BA: rddata <= 8'hE1; 14'h21BB: rddata <= 8'h30;
            14'h21BC: rddata <= 8'h02; 14'h21BD: rddata <= 8'hC5; 14'h21BE: rddata <= 8'hC9; 14'h21BF: rddata <= 8'hD6;
            14'h21C0: rddata <= 8'h54; 14'h21C1: rddata <= 8'hDA; 14'h21C2: rddata <= 8'hC4; 14'h21C3: rddata <= 8'h03;
            14'h21C4: rddata <= 8'hFE; 14'h21C5: rddata <= 8'h0D; 14'h21C6: rddata <= 8'hD2; 14'h21C7: rddata <= 8'hC4;
            14'h21C8: rddata <= 8'h03; 14'h21C9: rddata <= 8'h07; 14'h21CA: rddata <= 8'h4F; 14'h21CB: rddata <= 8'h06;
            14'h21CC: rddata <= 8'h00; 14'h21CD: rddata <= 8'hEB; 14'h21CE: rddata <= 8'h21; 14'h21CF: rddata <= 8'h5F;
            14'h21D0: rddata <= 8'h21; 14'h21D1: rddata <= 8'hC3; 14'h21D2: rddata <= 8'h65; 14'h21D3: rddata <= 8'h06;
            14'h21D4: rddata <= 8'hF1; 14'h21D5: rddata <= 8'hF1; 14'h21D6: rddata <= 8'hE1; 14'h21D7: rddata <= 8'hCA;
            14'h21D8: rddata <= 8'hCB; 14'h21D9: rddata <= 8'h0B; 14'h21DA: rddata <= 8'hE5; 14'h21DB: rddata <= 8'hCD;
            14'h21DC: rddata <= 8'h85; 14'h21DD: rddata <= 8'h09; 14'h21DE: rddata <= 8'hE1; 14'h21DF: rddata <= 8'h3A;
            14'h21E0: rddata <= 8'hAB; 14'h21E1: rddata <= 8'h38; 14'h21E2: rddata <= 8'h3D; 14'h21E3: rddata <= 8'hCA;
            14'h21E4: rddata <= 8'hA5; 14'h21E5: rddata <= 8'h28; 14'h21E6: rddata <= 8'hCD; 14'h21E7: rddata <= 8'hCF;
            14'h21E8: rddata <= 8'h0B; 14'h21E9: rddata <= 8'h01; 14'h21EA: rddata <= 8'h2C; 14'h21EB: rddata <= 8'h06;
            14'h21EC: rddata <= 8'hC3; 14'h21ED: rddata <= 8'hDB; 14'h21EE: rddata <= 8'h06; 14'h21EF: rddata <= 8'hC9;
            14'h21F0: rddata <= 8'h3E; 14'h21F1: rddata <= 8'h0B; 14'h21F2: rddata <= 8'hDF; 14'h21F3: rddata <= 8'hC9;
            14'h21F4: rddata <= 8'hCD; 14'h21F5: rddata <= 8'h72; 14'h21F6: rddata <= 8'h09; 14'h21F7: rddata <= 8'hCD;
            14'h21F8: rddata <= 8'h82; 14'h21F9: rddata <= 8'h06; 14'h21FA: rddata <= 8'hD5; 14'h21FB: rddata <= 8'hCF;
            14'h21FC: rddata <= 8'h2C; 14'h21FD: rddata <= 8'hCD; 14'h21FE: rddata <= 8'h54; 14'h21FF: rddata <= 8'h0B;
            14'h2200: rddata <= 8'hC1; 14'h2201: rddata <= 8'hED; 14'h2202: rddata <= 8'h79; 14'h2203: rddata <= 8'hC9;
            14'h2204: rddata <= 8'hCD; 14'h2205: rddata <= 8'h54; 14'h2206: rddata <= 8'h0B; 14'h2207: rddata <= 8'hF5;
            14'h2208: rddata <= 8'h3D; 14'h2209: rddata <= 8'hFE; 14'h220A: rddata <= 8'h26; 14'h220B: rddata <= 8'hD2;
            14'h220C: rddata <= 8'h97; 14'h220D: rddata <= 8'h06; 14'h220E: rddata <= 8'hCF; 14'h220F: rddata <= 8'h2C;
            14'h2210: rddata <= 8'hCD; 14'h2211: rddata <= 8'h54; 14'h2212: rddata <= 8'h0B; 14'h2213: rddata <= 8'hFE;
            14'h2214: rddata <= 8'h18; 14'h2215: rddata <= 8'hD2; 14'h2216: rddata <= 8'h97; 14'h2217: rddata <= 8'h06;
            14'h2218: rddata <= 8'h1C; 14'h2219: rddata <= 8'hF1; 14'h221A: rddata <= 8'h57; 14'h221B: rddata <= 8'hEB;
            14'h221C: rddata <= 8'hCD; 14'h221D: rddata <= 8'h21; 14'h221E: rddata <= 8'h22; 14'h221F: rddata <= 8'hEB;
            14'h2220: rddata <= 8'hC9; 14'h2221: rddata <= 8'hF5; 14'h2222: rddata <= 8'hE5; 14'h2223: rddata <= 8'hD9;
            14'h2224: rddata <= 8'h2A; 14'h2225: rddata <= 8'h01; 14'h2226: rddata <= 8'h38; 14'h2227: rddata <= 8'h3A;
            14'h2228: rddata <= 8'h0D; 14'h2229: rddata <= 8'h38; 14'h222A: rddata <= 8'h77; 14'h222B: rddata <= 8'hE1;
            14'h222C: rddata <= 8'h7D; 14'h222D: rddata <= 8'h87; 14'h222E: rddata <= 8'h87; 14'h222F: rddata <= 8'h85;
            14'h2230: rddata <= 8'hEB; 14'h2231: rddata <= 8'h5A; 14'h2232: rddata <= 8'h16; 14'h2233: rddata <= 8'h00;
            14'h2234: rddata <= 8'h62; 14'h2235: rddata <= 8'h6F; 14'h2236: rddata <= 8'h7B; 14'h2237: rddata <= 8'h3D;
            14'h2238: rddata <= 8'h29; 14'h2239: rddata <= 8'h29; 14'h223A: rddata <= 8'h29; 14'h223B: rddata <= 8'h19;
            14'h223C: rddata <= 8'h11; 14'h223D: rddata <= 8'h00; 14'h223E: rddata <= 8'h30; 14'h223F: rddata <= 8'h19;
            14'h2240: rddata <= 8'hC3; 14'h2241: rddata <= 8'hE7; 14'h2242: rddata <= 8'h1D; 14'h2243: rddata <= 8'hFE;
            14'h2244: rddata <= 8'h00; 14'h2245: rddata <= 8'hCA; 14'h2246: rddata <= 8'hD6; 14'h2247: rddata <= 8'h03;
            14'h2248: rddata <= 8'hCD; 14'h2249: rddata <= 8'h54; 14'h224A: rddata <= 8'h0B; 14'h224B: rddata <= 8'hFE;
            14'h224C: rddata <= 8'h10; 14'h224D: rddata <= 8'h30; 14'h224E: rddata <= 8'h10; 14'h224F: rddata <= 8'hD3;
            14'h2250: rddata <= 8'hF7; 14'h2251: rddata <= 8'hCF; 14'h2252: rddata <= 8'h2C; 14'h2253: rddata <= 8'hCD;
            14'h2254: rddata <= 8'h54; 14'h2255: rddata <= 8'h0B; 14'h2256: rddata <= 8'hD3; 14'h2257: rddata <= 8'hF6;
            14'h2258: rddata <= 8'h7E; 14'h2259: rddata <= 8'hFE; 14'h225A: rddata <= 8'h2C; 14'h225B: rddata <= 8'hC0;
            14'h225C: rddata <= 8'h23; 14'h225D: rddata <= 8'h18; 14'h225E: rddata <= 8'hE9; 14'h225F: rddata <= 8'hD6;
            14'h2260: rddata <= 8'h10; 14'h2261: rddata <= 8'hD3; 14'h2262: rddata <= 8'hF9; 14'h2263: rddata <= 8'hCF;
            14'h2264: rddata <= 8'h2C; 14'h2265: rddata <= 8'hCD; 14'h2266: rddata <= 8'h54; 14'h2267: rddata <= 8'h0B;
            14'h2268: rddata <= 8'hD3; 14'h2269: rddata <= 8'hF8; 14'h226A: rddata <= 8'h18; 14'h226B: rddata <= 8'hEC;
            14'h226C: rddata <= 8'hE1; 14'h226D: rddata <= 8'h23; 14'h226E: rddata <= 8'hCD; 14'h226F: rddata <= 8'h37;
            14'h2270: rddata <= 8'h0A; 14'h2271: rddata <= 8'hE3; 14'h2272: rddata <= 8'h11; 14'h2273: rddata <= 8'h49;
            14'h2274: rddata <= 8'h0A; 14'h2275: rddata <= 8'hD5; 14'h2276: rddata <= 8'hCD; 14'h2277: rddata <= 8'h82;
            14'h2278: rddata <= 8'h06; 14'h2279: rddata <= 8'h42; 14'h227A: rddata <= 8'h4B; 14'h227B: rddata <= 8'hED;
            14'h227C: rddata <= 8'h78; 14'h227D: rddata <= 8'hC3; 14'h227E: rddata <= 8'h36; 14'h227F: rddata <= 8'h0B;
            14'h2280: rddata <= 8'hE1; 14'h2281: rddata <= 8'h23; 14'h2282: rddata <= 8'hCD; 14'h2283: rddata <= 8'h37;
            14'h2284: rddata <= 8'h0A; 14'h2285: rddata <= 8'hE3; 14'h2286: rddata <= 8'h11; 14'h2287: rddata <= 8'h49;
            14'h2288: rddata <= 8'h0A; 14'h2289: rddata <= 8'hD5; 14'h228A: rddata <= 8'hCD; 14'h228B: rddata <= 8'h82;
            14'h228C: rddata <= 8'h06; 14'h228D: rddata <= 8'h7B; 14'h228E: rddata <= 8'hB7; 14'h228F: rddata <= 8'h20;
            14'h2290: rddata <= 8'h02; 14'h2291: rddata <= 8'h3E; 14'h2292: rddata <= 8'h03; 14'h2293: rddata <= 8'h5F;
            14'h2294: rddata <= 8'h01; 14'h2295: rddata <= 8'hF7; 14'h2296: rddata <= 8'h00; 14'h2297: rddata <= 8'h3E;
            14'h2298: rddata <= 8'hFF; 14'h2299: rddata <= 8'hCB; 14'h229A: rddata <= 8'h43; 14'h229B: rddata <= 8'h28;
            14'h229C: rddata <= 8'h0F; 14'h229D: rddata <= 8'h3E; 14'h229E: rddata <= 8'h0E; 14'h229F: rddata <= 8'hED;
            14'h22A0: rddata <= 8'h79; 14'h22A1: rddata <= 8'h0D; 14'h22A2: rddata <= 8'h06; 14'h22A3: rddata <= 8'hFF;
            14'h22A4: rddata <= 8'hED; 14'h22A5: rddata <= 8'h78; 14'h22A6: rddata <= 8'h10; 14'h22A7: rddata <= 8'hFC;
            14'h22A8: rddata <= 8'hFE; 14'h22A9: rddata <= 8'hFF; 14'h22AA: rddata <= 8'h20; 14'h22AB: rddata <= 8'h12;
            14'h22AC: rddata <= 8'hCB; 14'h22AD: rddata <= 8'h4B; 14'h22AE: rddata <= 8'h28; 14'h22AF: rddata <= 8'h0E;
            14'h22B0: rddata <= 8'h01; 14'h22B1: rddata <= 8'hF7; 14'h22B2: rddata <= 8'h00; 14'h22B3: rddata <= 8'h3E;
            14'h22B4: rddata <= 8'h0F; 14'h22B5: rddata <= 8'hED; 14'h22B6: rddata <= 8'h79; 14'h22B7: rddata <= 8'h0D;
            14'h22B8: rddata <= 8'h06; 14'h22B9: rddata <= 8'hFF; 14'h22BA: rddata <= 8'hED; 14'h22BB: rddata <= 8'h78;
            14'h22BC: rddata <= 8'h10; 14'h22BD: rddata <= 8'hFC; 14'h22BE: rddata <= 8'h2F; 14'h22BF: rddata <= 8'hC3;
            14'h22C0: rddata <= 8'h36; 14'h22C1: rddata <= 8'h0B; 14'h22C2: rddata <= 8'hE1; 14'h22C3: rddata <= 8'h23;
            14'h22C4: rddata <= 8'hCD; 14'h22C5: rddata <= 8'h37; 14'h22C6: rddata <= 8'h0A; 14'h22C7: rddata <= 8'hE3;
            14'h22C8: rddata <= 8'h11; 14'h22C9: rddata <= 8'h49; 14'h22CA: rddata <= 8'h0A; 14'h22CB: rddata <= 8'hD5;
            14'h22CC: rddata <= 8'hCD; 14'h22CD: rddata <= 8'h82; 14'h22CE: rddata <= 8'h06; 14'h22CF: rddata <= 8'h21;
            14'h22D0: rddata <= 8'hE9; 14'h22D1: rddata <= 8'h38; 14'h22D2: rddata <= 8'h7A; 14'h22D3: rddata <= 8'hB7;
            14'h22D4: rddata <= 8'h28; 14'h22D5: rddata <= 8'h04; 14'h22D6: rddata <= 8'h7A; 14'h22D7: rddata <= 8'hCD;
            14'h22D8: rddata <= 8'hE6; 14'h22D9: rddata <= 8'h22; 14'h22DA: rddata <= 8'h7B; 14'h22DB: rddata <= 8'hCD;
            14'h22DC: rddata <= 8'hE6; 14'h22DD: rddata <= 8'h22; 14'h22DE: rddata <= 8'h36; 14'h22DF: rddata <= 8'h00;
            14'h22E0: rddata <= 8'h21; 14'h22E1: rddata <= 8'hE9; 14'h22E2: rddata <= 8'h38; 14'h22E3: rddata <= 8'hC3;
            14'h22E4: rddata <= 8'h2F; 14'h22E5: rddata <= 8'h0E; 14'h22E6: rddata <= 8'h47; 14'h22E7: rddata <= 8'h1F;
            14'h22E8: rddata <= 8'h1F; 14'h22E9: rddata <= 8'h1F; 14'h22EA: rddata <= 8'h1F; 14'h22EB: rddata <= 8'hCD;
            14'h22EC: rddata <= 8'hEF; 14'h22ED: rddata <= 8'h22; 14'h22EE: rddata <= 8'h78; 14'h22EF: rddata <= 8'hE6;
            14'h22F0: rddata <= 8'h0F; 14'h22F1: rddata <= 8'hFE; 14'h22F2: rddata <= 8'h0A; 14'h22F3: rddata <= 8'h38;
            14'h22F4: rddata <= 8'h02; 14'h22F5: rddata <= 8'hC6; 14'h22F6: rddata <= 8'h07; 14'h22F7: rddata <= 8'hC6;
            14'h22F8: rddata <= 8'h30; 14'h22F9: rddata <= 8'h77; 14'h22FA: rddata <= 8'h23; 14'h22FB: rddata <= 8'hC9;
            14'h22FC: rddata <= 8'hCD; 14'h22FD: rddata <= 8'h72; 14'h22FE: rddata <= 8'h09; 14'h22FF: rddata <= 8'hCD;
            14'h2300: rddata <= 8'h82; 14'h2301: rddata <= 8'h06; 14'h2302: rddata <= 8'hD5; 14'h2303: rddata <= 8'hC9;
            14'h2304: rddata <= 8'hCD; 14'h2305: rddata <= 8'hE8; 14'h2306: rddata <= 8'h26; 14'h2307: rddata <= 8'hCD;
            14'h2308: rddata <= 8'hB4; 14'h2309: rddata <= 8'h26; 14'h230A: rddata <= 8'hCD; 14'h230B: rddata <= 8'h87;
            14'h230C: rddata <= 8'h27; 14'h230D: rddata <= 8'hFE; 14'h230E: rddata <= 8'h2C; 14'h230F: rddata <= 8'hC2;
            14'h2310: rddata <= 8'hF3; 14'h2311: rddata <= 8'h27; 14'h2312: rddata <= 8'hCD; 14'h2313: rddata <= 8'h86;
            14'h2314: rddata <= 8'h27; 14'h2315: rddata <= 8'hFE; 14'h2316: rddata <= 8'hAA; 14'h2317: rddata <= 8'h28;
            14'h2318: rddata <= 8'h0D; 14'h2319: rddata <= 8'hCD; 14'h231A: rddata <= 8'h72; 14'h231B: rddata <= 8'h09;
            14'h231C: rddata <= 8'hCD; 14'h231D: rddata <= 8'h82; 14'h231E: rddata <= 8'h06; 14'h231F: rddata <= 8'hED;
            14'h2320: rddata <= 8'h53; 14'h2321: rddata <= 8'hFC; 14'h2322: rddata <= 8'hBF; 14'h2323: rddata <= 8'hC3;
            14'h2324: rddata <= 8'hB3; 14'h2325: rddata <= 8'h27; 14'h2326: rddata <= 8'hCD; 14'h2327: rddata <= 8'h2C;
            14'h2328: rddata <= 8'h23; 14'h2329: rddata <= 8'hC3; 14'h232A: rddata <= 8'hC5; 14'h232B: rddata <= 8'h27;
            14'h232C: rddata <= 8'h23; 14'h232D: rddata <= 8'h3E; 14'h232E: rddata <= 8'h01; 14'h232F: rddata <= 8'h32;
            14'h2330: rddata <= 8'hCB; 14'h2331: rddata <= 8'h38; 14'h2332: rddata <= 8'hCD; 14'h2333: rddata <= 8'hD1;
            14'h2334: rddata <= 8'h10; 14'h2335: rddata <= 8'h32; 14'h2336: rddata <= 8'hCB; 14'h2337: rddata <= 8'h38;
            14'h2338: rddata <= 8'hC2; 14'h2339: rddata <= 8'h97; 14'h233A: rddata <= 8'h06; 14'h233B: rddata <= 8'hCD;
            14'h233C: rddata <= 8'h75; 14'h233D: rddata <= 8'h09; 14'h233E: rddata <= 8'hE5; 14'h233F: rddata <= 8'h60;
            14'h2340: rddata <= 8'h69; 14'h2341: rddata <= 8'h4E; 14'h2342: rddata <= 8'h06; 14'h2343: rddata <= 8'h00;
            14'h2344: rddata <= 8'h09; 14'h2345: rddata <= 8'h09; 14'h2346: rddata <= 8'h23; 14'h2347: rddata <= 8'h22;
            14'h2348: rddata <= 8'hFC; 14'h2349: rddata <= 8'hBF; 14'h234A: rddata <= 8'h1B; 14'h234B: rddata <= 8'h1B;
            14'h234C: rddata <= 8'h1B; 14'h234D: rddata <= 8'hED; 14'h234E: rddata <= 8'h53; 14'h234F: rddata <= 8'hFE;
            14'h2350: rddata <= 8'hBF; 14'h2351: rddata <= 8'hE1; 14'h2352: rddata <= 8'hC9; 14'h2353: rddata <= 8'hCD;
            14'h2354: rddata <= 8'hE8; 14'h2355: rddata <= 8'h26; 14'h2356: rddata <= 8'hCD; 14'h2357: rddata <= 8'hB4;
            14'h2358: rddata <= 8'h26; 14'h2359: rddata <= 8'hCD; 14'h235A: rddata <= 8'h87; 14'h235B: rddata <= 8'h27;
            14'h235C: rddata <= 8'hFE; 14'h235D: rddata <= 8'h2C; 14'h235E: rddata <= 8'hC2; 14'h235F: rddata <= 8'h30;
            14'h2360: rddata <= 8'h28; 14'h2361: rddata <= 8'hCD; 14'h2362: rddata <= 8'h86; 14'h2363: rddata <= 8'h27;
            14'h2364: rddata <= 8'hFE; 14'h2365: rddata <= 8'hAA; 14'h2366: rddata <= 8'h28; 14'h2367: rddata <= 8'h20;
            14'h2368: rddata <= 8'hCD; 14'h2369: rddata <= 8'h72; 14'h236A: rddata <= 8'h09; 14'h236B: rddata <= 8'hCD;
            14'h236C: rddata <= 8'h82; 14'h236D: rddata <= 8'h06; 14'h236E: rddata <= 8'hED; 14'h236F: rddata <= 8'h53;
            14'h2370: rddata <= 8'hFC; 14'h2371: rddata <= 8'hBF; 14'h2372: rddata <= 8'hCD; 14'h2373: rddata <= 8'h87;
            14'h2374: rddata <= 8'h27; 14'h2375: rddata <= 8'hFE; 14'h2376: rddata <= 8'h2C; 14'h2377: rddata <= 8'hC2;
            14'h2378: rddata <= 8'hD6; 14'h2379: rddata <= 8'h03; 14'h237A: rddata <= 8'h23; 14'h237B: rddata <= 8'hCD;
            14'h237C: rddata <= 8'h72; 14'h237D: rddata <= 8'h09; 14'h237E: rddata <= 8'hCD; 14'h237F: rddata <= 8'h82;
            14'h2380: rddata <= 8'h06; 14'h2381: rddata <= 8'hED; 14'h2382: rddata <= 8'h53; 14'h2383: rddata <= 8'hFE;
            14'h2384: rddata <= 8'hBF; 14'h2385: rddata <= 8'hC3; 14'h2386: rddata <= 8'h92; 14'h2387: rddata <= 8'h28;
            14'h2388: rddata <= 8'hCD; 14'h2389: rddata <= 8'h2C; 14'h238A: rddata <= 8'h23; 14'h238B: rddata <= 8'hC3;
            14'h238C: rddata <= 8'h67; 14'h238D: rddata <= 8'h28; 14'h238E: rddata <= 8'hCD; 14'h238F: rddata <= 8'hB4;
            14'h2390: rddata <= 8'h26; 14'h2391: rddata <= 8'hE5; 14'h2392: rddata <= 8'h3E; 14'h2393: rddata <= 8'h19;
            14'h2394: rddata <= 8'hCD; 14'h2395: rddata <= 8'hEF; 14'h2396: rddata <= 8'h25; 14'h2397: rddata <= 8'hCD;
            14'h2398: rddata <= 8'hD3; 14'h2399: rddata <= 8'h26; 14'h239A: rddata <= 8'hCD; 14'h239B: rddata <= 8'hE0;
            14'h239C: rddata <= 8'h26; 14'h239D: rddata <= 8'hE1; 14'h239E: rddata <= 8'hC9; 14'h239F: rddata <= 8'hE5;
            14'h23A0: rddata <= 8'hB7; 14'h23A1: rddata <= 8'h20; 14'h23A2: rddata <= 8'h18; 14'h23A3: rddata <= 8'h3E;
            14'h23A4: rddata <= 8'h1E; 14'h23A5: rddata <= 8'hCD; 14'h23A6: rddata <= 8'hEF; 14'h23A7: rddata <= 8'h25;
            14'h23A8: rddata <= 8'hCD; 14'h23A9: rddata <= 8'hE0; 14'h23AA: rddata <= 8'h26; 14'h23AB: rddata <= 8'hCD;
            14'h23AC: rddata <= 8'h02; 14'h23AD: rddata <= 8'h26; 14'h23AE: rddata <= 8'hB7; 14'h23AF: rddata <= 8'h28;
            14'h23B0: rddata <= 8'h05; 14'h23B1: rddata <= 8'hCD; 14'h23B2: rddata <= 8'h72; 14'h23B3: rddata <= 8'h1D;
            14'h23B4: rddata <= 8'h18; 14'h23B5: rddata <= 8'hF5; 14'h23B6: rddata <= 8'hCD; 14'h23B7: rddata <= 8'hEA;
            14'h23B8: rddata <= 8'h19; 14'h23B9: rddata <= 8'hE1; 14'h23BA: rddata <= 8'hC9; 14'h23BB: rddata <= 8'hE1;
            14'h23BC: rddata <= 8'hCD; 14'h23BD: rddata <= 8'hB4; 14'h23BE: rddata <= 8'h26; 14'h23BF: rddata <= 8'hE5;
            14'h23C0: rddata <= 8'h3E; 14'h23C1: rddata <= 8'h1C; 14'h23C2: rddata <= 8'hCD; 14'h23C3: rddata <= 8'hEF;
            14'h23C4: rddata <= 8'h25; 14'h23C5: rddata <= 8'hCD; 14'h23C6: rddata <= 8'hD3; 14'h23C7: rddata <= 8'h26;
            14'h23C8: rddata <= 8'hCD; 14'h23C9: rddata <= 8'hE0; 14'h23CA: rddata <= 8'h26; 14'h23CB: rddata <= 8'h18;
            14'h23CC: rddata <= 8'hEC; 14'h23CD: rddata <= 8'hCD; 14'h23CE: rddata <= 8'hB4; 14'h23CF: rddata <= 8'h26;
            14'h23D0: rddata <= 8'hE5; 14'h23D1: rddata <= 8'h3E; 14'h23D2: rddata <= 8'h1B; 14'h23D3: rddata <= 8'hCD;
            14'h23D4: rddata <= 8'hEF; 14'h23D5: rddata <= 8'h25; 14'h23D6: rddata <= 8'hCD; 14'h23D7: rddata <= 8'hD3;
            14'h23D8: rddata <= 8'h26; 14'h23D9: rddata <= 8'hCD; 14'h23DA: rddata <= 8'hE0; 14'h23DB: rddata <= 8'h26;
            14'h23DC: rddata <= 8'hE1; 14'h23DD: rddata <= 8'hC9; 14'h23DE: rddata <= 8'hE5; 14'h23DF: rddata <= 8'hB7;
            14'h23E0: rddata <= 8'h20; 14'h23E1: rddata <= 8'h09; 14'h23E2: rddata <= 8'hAF; 14'h23E3: rddata <= 8'h32;
            14'h23E4: rddata <= 8'h00; 14'h23E5: rddata <= 8'hBF; 14'h23E6: rddata <= 8'h32; 14'h23E7: rddata <= 8'h01;
            14'h23E8: rddata <= 8'hBF; 14'h23E9: rddata <= 8'h18; 14'h23EA: rddata <= 8'h05; 14'h23EB: rddata <= 8'hE1;
            14'h23EC: rddata <= 8'hCD; 14'h23ED: rddata <= 8'hB4; 14'h23EE: rddata <= 8'h26; 14'h23EF: rddata <= 8'hE5;
            14'h23F0: rddata <= 8'hCD; 14'h23F1: rddata <= 8'hE8; 14'h23F2: rddata <= 8'h26; 14'h23F3: rddata <= 8'h3E;
            14'h23F4: rddata <= 8'h16; 14'h23F5: rddata <= 8'hCD; 14'h23F6: rddata <= 8'hEF; 14'h23F7: rddata <= 8'h25;
            14'h23F8: rddata <= 8'hCD; 14'h23F9: rddata <= 8'hD3; 14'h23FA: rddata <= 8'h26; 14'h23FB: rddata <= 8'hCD;
            14'h23FC: rddata <= 8'hE0; 14'h23FD: rddata <= 8'h26; 14'h23FE: rddata <= 8'h3E; 14'h23FF: rddata <= 8'h18;
            14'h2400: rddata <= 8'h32; 14'h2401: rddata <= 8'h08; 14'h2402: rddata <= 8'h38; 14'h2403: rddata <= 8'h3E;
            14'h2404: rddata <= 8'h18; 14'h2405: rddata <= 8'hCD; 14'h2406: rddata <= 8'hEF; 14'h2407: rddata <= 8'h25;
            14'h2408: rddata <= 8'hAF; 14'h2409: rddata <= 8'hCD; 14'h240A: rddata <= 8'h0B; 14'h240B: rddata <= 8'h26;
            14'h240C: rddata <= 8'hCD; 14'h240D: rddata <= 8'h02; 14'h240E: rddata <= 8'h26; 14'h240F: rddata <= 8'hFE;
            14'h2410: rddata <= 8'hFC; 14'h2411: rddata <= 8'hCA; 14'h2412: rddata <= 8'h45; 14'h2413: rddata <= 8'h25;
            14'h2414: rddata <= 8'hB7; 14'h2415: rddata <= 8'hF2; 14'h2416: rddata <= 8'h1C; 14'h2417: rddata <= 8'h24;
            14'h2418: rddata <= 8'hE1; 14'h2419: rddata <= 8'hC3; 14'h241A: rddata <= 8'h57; 14'h241B: rddata <= 8'h25;
            14'h241C: rddata <= 8'hCD; 14'h241D: rddata <= 8'h02; 14'h241E: rddata <= 8'h26; 14'h241F: rddata <= 8'h32;
            14'h2420: rddata <= 8'h52; 14'h2421: rddata <= 8'h38; 14'h2422: rddata <= 8'hCD; 14'h2423: rddata <= 8'h02;
            14'h2424: rddata <= 8'h26; 14'h2425: rddata <= 8'h32; 14'h2426: rddata <= 8'h53; 14'h2427: rddata <= 8'h38;
            14'h2428: rddata <= 8'hCB; 14'h2429: rddata <= 8'h3F; 14'h242A: rddata <= 8'hC6; 14'h242B: rddata <= 8'h50;
            14'h242C: rddata <= 8'hCD; 14'h242D: rddata <= 8'h16; 14'h242E: rddata <= 8'h26; 14'h242F: rddata <= 8'h3E;
            14'h2430: rddata <= 8'h2D; 14'h2431: rddata <= 8'hCD; 14'h2432: rddata <= 8'h72; 14'h2433: rddata <= 8'h1D;
            14'h2434: rddata <= 8'h3A; 14'h2435: rddata <= 8'h53; 14'h2436: rddata <= 8'h38; 14'h2437: rddata <= 8'h1F;
            14'h2438: rddata <= 8'h3A; 14'h2439: rddata <= 8'h52; 14'h243A: rddata <= 8'h38; 14'h243B: rddata <= 8'h1F;
            14'h243C: rddata <= 8'hCB; 14'h243D: rddata <= 8'h3F; 14'h243E: rddata <= 8'hCB; 14'h243F: rddata <= 8'h3F;
            14'h2440: rddata <= 8'hCB; 14'h2441: rddata <= 8'h3F; 14'h2442: rddata <= 8'hCB; 14'h2443: rddata <= 8'h3F;
            14'h2444: rddata <= 8'hCD; 14'h2445: rddata <= 8'h16; 14'h2446: rddata <= 8'h26; 14'h2447: rddata <= 8'h3E;
            14'h2448: rddata <= 8'h2D; 14'h2449: rddata <= 8'hCD; 14'h244A: rddata <= 8'h72; 14'h244B: rddata <= 8'h1D;
            14'h244C: rddata <= 8'h3A; 14'h244D: rddata <= 8'h52; 14'h244E: rddata <= 8'h38; 14'h244F: rddata <= 8'hE6;
            14'h2450: rddata <= 8'h1F; 14'h2451: rddata <= 8'hCD; 14'h2452: rddata <= 8'h16; 14'h2453: rddata <= 8'h26;
            14'h2454: rddata <= 8'h3E; 14'h2455: rddata <= 8'h20; 14'h2456: rddata <= 8'hCD; 14'h2457: rddata <= 8'h72;
            14'h2458: rddata <= 8'h1D; 14'h2459: rddata <= 8'hCD; 14'h245A: rddata <= 8'h02; 14'h245B: rddata <= 8'h26;
            14'h245C: rddata <= 8'h32; 14'h245D: rddata <= 8'h52; 14'h245E: rddata <= 8'h38; 14'h245F: rddata <= 8'hCD;
            14'h2460: rddata <= 8'h02; 14'h2461: rddata <= 8'h26; 14'h2462: rddata <= 8'h32; 14'h2463: rddata <= 8'h53;
            14'h2464: rddata <= 8'h38; 14'h2465: rddata <= 8'hCB; 14'h2466: rddata <= 8'h3F; 14'h2467: rddata <= 8'hCB;
            14'h2468: rddata <= 8'h3F; 14'h2469: rddata <= 8'hCB; 14'h246A: rddata <= 8'h3F; 14'h246B: rddata <= 8'hCD;
            14'h246C: rddata <= 8'h16; 14'h246D: rddata <= 8'h26; 14'h246E: rddata <= 8'h3E; 14'h246F: rddata <= 8'h3A;
            14'h2470: rddata <= 8'hCD; 14'h2471: rddata <= 8'h72; 14'h2472: rddata <= 8'h1D; 14'h2473: rddata <= 8'h3A;
            14'h2474: rddata <= 8'h53; 14'h2475: rddata <= 8'h38; 14'h2476: rddata <= 8'hE6; 14'h2477: rddata <= 8'h07;
            14'h2478: rddata <= 8'h4F; 14'h2479: rddata <= 8'h3A; 14'h247A: rddata <= 8'h52; 14'h247B: rddata <= 8'h38;
            14'h247C: rddata <= 8'hCB; 14'h247D: rddata <= 8'h39; 14'h247E: rddata <= 8'h1F; 14'h247F: rddata <= 8'hCB;
            14'h2480: rddata <= 8'h39; 14'h2481: rddata <= 8'h1F; 14'h2482: rddata <= 8'hCB; 14'h2483: rddata <= 8'h39;
            14'h2484: rddata <= 8'h1F; 14'h2485: rddata <= 8'hCB; 14'h2486: rddata <= 8'h39; 14'h2487: rddata <= 8'h1F;
            14'h2488: rddata <= 8'hCB; 14'h2489: rddata <= 8'h39; 14'h248A: rddata <= 8'h1F; 14'h248B: rddata <= 8'hCD;
            14'h248C: rddata <= 8'h16; 14'h248D: rddata <= 8'h26; 14'h248E: rddata <= 8'hCD; 14'h248F: rddata <= 8'h02;
            14'h2490: rddata <= 8'h26; 14'h2491: rddata <= 8'hCB; 14'h2492: rddata <= 8'h47; 14'h2493: rddata <= 8'h28;
            14'h2494: rddata <= 8'h14; 14'h2495: rddata <= 8'h21; 14'h2496: rddata <= 8'h3E; 14'h2497: rddata <= 8'h25;
            14'h2498: rddata <= 8'hCD; 14'h2499: rddata <= 8'h9D; 14'h249A: rddata <= 8'h0E; 14'h249B: rddata <= 8'hCD;
            14'h249C: rddata <= 8'h02; 14'h249D: rddata <= 8'h26; 14'h249E: rddata <= 8'hCD; 14'h249F: rddata <= 8'h02;
            14'h24A0: rddata <= 8'h26; 14'h24A1: rddata <= 8'hCD; 14'h24A2: rddata <= 8'h02; 14'h24A3: rddata <= 8'h26;
            14'h24A4: rddata <= 8'hCD; 14'h24A5: rddata <= 8'h02; 14'h24A6: rddata <= 8'h26; 14'h24A7: rddata <= 8'h18;
            14'h24A8: rddata <= 8'h7F; 14'h24A9: rddata <= 8'hCD; 14'h24AA: rddata <= 8'h02; 14'h24AB: rddata <= 8'h26;
            14'h24AC: rddata <= 8'h32; 14'h24AD: rddata <= 8'h52; 14'h24AE: rddata <= 8'h38; 14'h24AF: rddata <= 8'hCD;
            14'h24B0: rddata <= 8'h02; 14'h24B1: rddata <= 8'h26; 14'h24B2: rddata <= 8'h32; 14'h24B3: rddata <= 8'h53;
            14'h24B4: rddata <= 8'h38; 14'h24B5: rddata <= 8'hCD; 14'h24B6: rddata <= 8'h02; 14'h24B7: rddata <= 8'h26;
            14'h24B8: rddata <= 8'h32; 14'h24B9: rddata <= 8'h54; 14'h24BA: rddata <= 8'h38; 14'h24BB: rddata <= 8'hCD;
            14'h24BC: rddata <= 8'h02; 14'h24BD: rddata <= 8'h26; 14'h24BE: rddata <= 8'h32; 14'h24BF: rddata <= 8'h55;
            14'h24C0: rddata <= 8'h38; 14'h24C1: rddata <= 8'hB7; 14'h24C2: rddata <= 8'h20; 14'h24C3: rddata <= 8'h42;
            14'h24C4: rddata <= 8'h3A; 14'h24C5: rddata <= 8'h54; 14'h24C6: rddata <= 8'h38; 14'h24C7: rddata <= 8'hE6;
            14'h24C8: rddata <= 8'hF0; 14'h24C9: rddata <= 8'h20; 14'h24CA: rddata <= 8'h3B; 14'h24CB: rddata <= 8'h3A;
            14'h24CC: rddata <= 8'h54; 14'h24CD: rddata <= 8'h38; 14'h24CE: rddata <= 8'hB7; 14'h24CF: rddata <= 8'h20;
            14'h24D0: rddata <= 8'h19; 14'h24D1: rddata <= 8'h3A; 14'h24D2: rddata <= 8'h53; 14'h24D3: rddata <= 8'h38;
            14'h24D4: rddata <= 8'hE6; 14'h24D5: rddata <= 8'hFC; 14'h24D6: rddata <= 8'h20; 14'h24D7: rddata <= 8'h12;
            14'h24D8: rddata <= 8'h3A; 14'h24D9: rddata <= 8'h53; 14'h24DA: rddata <= 8'h38; 14'h24DB: rddata <= 8'h67;
            14'h24DC: rddata <= 8'h3A; 14'h24DD: rddata <= 8'h52; 14'h24DE: rddata <= 8'h38; 14'h24DF: rddata <= 8'h6F;
            14'h24E0: rddata <= 8'hCD; 14'h24E1: rddata <= 8'h35; 14'h24E2: rddata <= 8'h26; 14'h24E3: rddata <= 8'h3E;
            14'h24E4: rddata <= 8'h42; 14'h24E5: rddata <= 8'hCD; 14'h24E6: rddata <= 8'h72; 14'h24E7: rddata <= 8'h1D;
            14'h24E8: rddata <= 8'h18; 14'h24E9: rddata <= 8'h3E; 14'h24EA: rddata <= 8'h3A; 14'h24EB: rddata <= 8'h54;
            14'h24EC: rddata <= 8'h38; 14'h24ED: rddata <= 8'hE6; 14'h24EE: rddata <= 8'h0F; 14'h24EF: rddata <= 8'h67;
            14'h24F0: rddata <= 8'h3A; 14'h24F1: rddata <= 8'h53; 14'h24F2: rddata <= 8'h38; 14'h24F3: rddata <= 8'h6F;
            14'h24F4: rddata <= 8'hCB; 14'h24F5: rddata <= 8'h3C; 14'h24F6: rddata <= 8'hCB; 14'h24F7: rddata <= 8'h1D;
            14'h24F8: rddata <= 8'hCB; 14'h24F9: rddata <= 8'h3C; 14'h24FA: rddata <= 8'hCB; 14'h24FB: rddata <= 8'h1D;
            14'h24FC: rddata <= 8'hCD; 14'h24FD: rddata <= 8'h35; 14'h24FE: rddata <= 8'h26; 14'h24FF: rddata <= 8'h3E;
            14'h2500: rddata <= 8'h4B; 14'h2501: rddata <= 8'hCD; 14'h2502: rddata <= 8'h72; 14'h2503: rddata <= 8'h1D;
            14'h2504: rddata <= 8'h18; 14'h2505: rddata <= 8'h22; 14'h2506: rddata <= 8'h3A; 14'h2507: rddata <= 8'h55;
            14'h2508: rddata <= 8'h38; 14'h2509: rddata <= 8'h67; 14'h250A: rddata <= 8'h3A; 14'h250B: rddata <= 8'h54;
            14'h250C: rddata <= 8'h38; 14'h250D: rddata <= 8'h6F; 14'h250E: rddata <= 8'hCB; 14'h250F: rddata <= 8'h3C;
            14'h2510: rddata <= 8'hCB; 14'h2511: rddata <= 8'h1D; 14'h2512: rddata <= 8'hCB; 14'h2513: rddata <= 8'h3C;
            14'h2514: rddata <= 8'hCB; 14'h2515: rddata <= 8'h1D; 14'h2516: rddata <= 8'hCB; 14'h2517: rddata <= 8'h3C;
            14'h2518: rddata <= 8'hCB; 14'h2519: rddata <= 8'h1D; 14'h251A: rddata <= 8'hCB; 14'h251B: rddata <= 8'h3C;
            14'h251C: rddata <= 8'hCB; 14'h251D: rddata <= 8'h1D; 14'h251E: rddata <= 8'hCD; 14'h251F: rddata <= 8'h35;
            14'h2520: rddata <= 8'h26; 14'h2521: rddata <= 8'h3E; 14'h2522: rddata <= 8'h4D; 14'h2523: rddata <= 8'hCD;
            14'h2524: rddata <= 8'h72; 14'h2525: rddata <= 8'h1D; 14'h2526: rddata <= 8'h18; 14'h2527: rddata <= 8'h00;
            14'h2528: rddata <= 8'h3E; 14'h2529: rddata <= 8'h20; 14'h252A: rddata <= 8'hCD; 14'h252B: rddata <= 8'h72;
            14'h252C: rddata <= 8'h1D; 14'h252D: rddata <= 8'hCD; 14'h252E: rddata <= 8'h02; 14'h252F: rddata <= 8'h26;
            14'h2530: rddata <= 8'hB7; 14'h2531: rddata <= 8'h28; 14'h2532: rddata <= 8'h05; 14'h2533: rddata <= 8'hCD;
            14'h2534: rddata <= 8'h72; 14'h2535: rddata <= 8'h1D; 14'h2536: rddata <= 8'h18; 14'h2537: rddata <= 8'hF5;
            14'h2538: rddata <= 8'hCD; 14'h2539: rddata <= 8'hEA; 14'h253A: rddata <= 8'h19; 14'h253B: rddata <= 8'hC3;
            14'h253C: rddata <= 8'h03; 14'h253D: rddata <= 8'h24; 14'h253E: rddata <= 8'h20; 14'h253F: rddata <= 8'h3C;
            14'h2540: rddata <= 8'h44; 14'h2541: rddata <= 8'h49; 14'h2542: rddata <= 8'h52; 14'h2543: rddata <= 8'h3E;
            14'h2544: rddata <= 8'h00; 14'h2545: rddata <= 8'h3E; 14'h2546: rddata <= 8'h17; 14'h2547: rddata <= 8'hCD;
            14'h2548: rddata <= 8'hEF; 14'h2549: rddata <= 8'h25; 14'h254A: rddata <= 8'hAF; 14'h254B: rddata <= 8'hCD;
            14'h254C: rddata <= 8'h0B; 14'h254D: rddata <= 8'h26; 14'h254E: rddata <= 8'hCD; 14'h254F: rddata <= 8'h02;
            14'h2550: rddata <= 8'h26; 14'h2551: rddata <= 8'hB7; 14'h2552: rddata <= 8'hFA; 14'h2553: rddata <= 8'h57;
            14'h2554: rddata <= 8'h25; 14'h2555: rddata <= 8'hE1; 14'h2556: rddata <= 8'hC9; 14'h2557: rddata <= 8'hED;
            14'h2558: rddata <= 8'h44; 14'h2559: rddata <= 8'h3D; 14'h255A: rddata <= 8'hFE; 14'h255B: rddata <= 8'h08;
            14'h255C: rddata <= 8'h38; 14'h255D: rddata <= 8'h02; 14'h255E: rddata <= 8'h3E; 14'h255F: rddata <= 8'h05;
            14'h2560: rddata <= 8'h21; 14'h2561: rddata <= 8'h74; 14'h2562: rddata <= 8'h25; 14'h2563: rddata <= 8'h87;
            14'h2564: rddata <= 8'h85; 14'h2565: rddata <= 8'h6F; 14'h2566: rddata <= 8'h7C; 14'h2567: rddata <= 8'hCE;
            14'h2568: rddata <= 8'h00; 14'h2569: rddata <= 8'h67; 14'h256A: rddata <= 8'h7E; 14'h256B: rddata <= 8'h23;
            14'h256C: rddata <= 8'h66; 14'h256D: rddata <= 8'h6F; 14'h256E: rddata <= 8'h3E; 14'h256F: rddata <= 8'h3F;
            14'h2570: rddata <= 8'hDF; 14'h2571: rddata <= 8'hC3; 14'h2572: rddata <= 8'hF4; 14'h2573: rddata <= 8'h03;
            14'h2574: rddata <= 8'h84; 14'h2575: rddata <= 8'h25; 14'h2576: rddata <= 8'h8E; 14'h2577: rddata <= 8'h25;
            14'h2578: rddata <= 8'h9C; 14'h2579: rddata <= 8'h25; 14'h257A: rddata <= 8'hAA; 14'h257B: rddata <= 8'h25;
            14'h257C: rddata <= 8'hAE; 14'h257D: rddata <= 8'h25; 14'h257E: rddata <= 8'hBD; 14'h257F: rddata <= 8'h25;
            14'h2580: rddata <= 8'hCB; 14'h2581: rddata <= 8'h25; 14'h2582: rddata <= 8'hD3; 14'h2583: rddata <= 8'h25;
            14'h2584: rddata <= 8'h4E; 14'h2585: rddata <= 8'h6F; 14'h2586: rddata <= 8'h74; 14'h2587: rddata <= 8'h20;
            14'h2588: rddata <= 8'h66; 14'h2589: rddata <= 8'h6F; 14'h258A: rddata <= 8'h75; 14'h258B: rddata <= 8'h6E;
            14'h258C: rddata <= 8'h64; 14'h258D: rddata <= 8'h00; 14'h258E: rddata <= 8'h54; 14'h258F: rddata <= 8'h6F;
            14'h2590: rddata <= 8'h6F; 14'h2591: rddata <= 8'h20; 14'h2592: rddata <= 8'h6D; 14'h2593: rddata <= 8'h61;
            14'h2594: rddata <= 8'h6E; 14'h2595: rddata <= 8'h79; 14'h2596: rddata <= 8'h20; 14'h2597: rddata <= 8'h6F;
            14'h2598: rddata <= 8'h70; 14'h2599: rddata <= 8'h65; 14'h259A: rddata <= 8'h6E; 14'h259B: rddata <= 8'h00;
            14'h259C: rddata <= 8'h49; 14'h259D: rddata <= 8'h6E; 14'h259E: rddata <= 8'h76; 14'h259F: rddata <= 8'h61;
            14'h25A0: rddata <= 8'h6C; 14'h25A1: rddata <= 8'h69; 14'h25A2: rddata <= 8'h64; 14'h25A3: rddata <= 8'h20;
            14'h25A4: rddata <= 8'h70; 14'h25A5: rddata <= 8'h61; 14'h25A6: rddata <= 8'h72; 14'h25A7: rddata <= 8'h61;
            14'h25A8: rddata <= 8'h6D; 14'h25A9: rddata <= 8'h00; 14'h25AA: rddata <= 8'h45; 14'h25AB: rddata <= 8'h4F;
            14'h25AC: rddata <= 8'h46; 14'h25AD: rddata <= 8'h00; 14'h25AE: rddata <= 8'h41; 14'h25AF: rddata <= 8'h6C;
            14'h25B0: rddata <= 8'h72; 14'h25B1: rddata <= 8'h65; 14'h25B2: rddata <= 8'h61; 14'h25B3: rddata <= 8'h64;
            14'h25B4: rddata <= 8'h79; 14'h25B5: rddata <= 8'h20; 14'h25B6: rddata <= 8'h65; 14'h25B7: rddata <= 8'h78;
            14'h25B8: rddata <= 8'h69; 14'h25B9: rddata <= 8'h73; 14'h25BA: rddata <= 8'h74; 14'h25BB: rddata <= 8'h73;
            14'h25BC: rddata <= 8'h00; 14'h25BD: rddata <= 8'h55; 14'h25BE: rddata <= 8'h6E; 14'h25BF: rddata <= 8'h6B;
            14'h25C0: rddata <= 8'h6E; 14'h25C1: rddata <= 8'h6F; 14'h25C2: rddata <= 8'h77; 14'h25C3: rddata <= 8'h6E;
            14'h25C4: rddata <= 8'h20; 14'h25C5: rddata <= 8'h65; 14'h25C6: rddata <= 8'h72; 14'h25C7: rddata <= 8'h72;
            14'h25C8: rddata <= 8'h6F; 14'h25C9: rddata <= 8'h72; 14'h25CA: rddata <= 8'h00; 14'h25CB: rddata <= 8'h4E;
            14'h25CC: rddata <= 8'h6F; 14'h25CD: rddata <= 8'h20; 14'h25CE: rddata <= 8'h64; 14'h25CF: rddata <= 8'h69;
            14'h25D0: rddata <= 8'h73; 14'h25D1: rddata <= 8'h6B; 14'h25D2: rddata <= 8'h00; 14'h25D3: rddata <= 8'h4E;
            14'h25D4: rddata <= 8'h6F; 14'h25D5: rddata <= 8'h74; 14'h25D6: rddata <= 8'h20; 14'h25D7: rddata <= 8'h65;
            14'h25D8: rddata <= 8'h6D; 14'h25D9: rddata <= 8'h70; 14'h25DA: rddata <= 8'h74; 14'h25DB: rddata <= 8'h79;
            14'h25DC: rddata <= 8'h00; 14'h25DD: rddata <= 8'h21; 14'h25DE: rddata <= 8'hE6; 14'h25DF: rddata <= 8'h25;
            14'h25E0: rddata <= 8'h3E; 14'h25E1: rddata <= 8'h3F; 14'h25E2: rddata <= 8'hDF; 14'h25E3: rddata <= 8'hC3;
            14'h25E4: rddata <= 8'hF4; 14'h25E5: rddata <= 8'h03; 14'h25E6: rddata <= 8'h42; 14'h25E7: rddata <= 8'h61;
            14'h25E8: rddata <= 8'h64; 14'h25E9: rddata <= 8'h20; 14'h25EA: rddata <= 8'h66; 14'h25EB: rddata <= 8'h69;
            14'h25EC: rddata <= 8'h6C; 14'h25ED: rddata <= 8'h65; 14'h25EE: rddata <= 8'h00; 14'h25EF: rddata <= 8'hF5;
            14'h25F0: rddata <= 8'hDB; 14'h25F1: rddata <= 8'hF4; 14'h25F2: rddata <= 8'hE6; 14'h25F3: rddata <= 8'h01;
            14'h25F4: rddata <= 8'h28; 14'h25F5: rddata <= 8'h04; 14'h25F6: rddata <= 8'hDB; 14'h25F7: rddata <= 8'hF5;
            14'h25F8: rddata <= 8'h18; 14'h25F9: rddata <= 8'hF6; 14'h25FA: rddata <= 8'h3E; 14'h25FB: rddata <= 8'h80;
            14'h25FC: rddata <= 8'hD3; 14'h25FD: rddata <= 8'hF4; 14'h25FE: rddata <= 8'hF1; 14'h25FF: rddata <= 8'hC3;
            14'h2600: rddata <= 8'h0B; 14'h2601: rddata <= 8'h26; 14'h2602: rddata <= 8'hDB; 14'h2603: rddata <= 8'hF4;
            14'h2604: rddata <= 8'hE6; 14'h2605: rddata <= 8'h01; 14'h2606: rddata <= 8'h28; 14'h2607: rddata <= 8'hFA;
            14'h2608: rddata <= 8'hDB; 14'h2609: rddata <= 8'hF5; 14'h260A: rddata <= 8'hC9; 14'h260B: rddata <= 8'hF5;
            14'h260C: rddata <= 8'hDB; 14'h260D: rddata <= 8'hF4; 14'h260E: rddata <= 8'hE6; 14'h260F: rddata <= 8'h02;
            14'h2610: rddata <= 8'h20; 14'h2611: rddata <= 8'hFA; 14'h2612: rddata <= 8'hF1; 14'h2613: rddata <= 8'hD3;
            14'h2614: rddata <= 8'hF5; 14'h2615: rddata <= 8'hC9; 14'h2616: rddata <= 8'hFE; 14'h2617: rddata <= 8'h64;
            14'h2618: rddata <= 8'h38; 14'h2619: rddata <= 8'h04; 14'h261A: rddata <= 8'hD6; 14'h261B: rddata <= 8'h64;
            14'h261C: rddata <= 8'h18; 14'h261D: rddata <= 8'hF8; 14'h261E: rddata <= 8'h0E; 14'h261F: rddata <= 8'h00;
            14'h2620: rddata <= 8'h0C; 14'h2621: rddata <= 8'hD6; 14'h2622: rddata <= 8'h0A; 14'h2623: rddata <= 8'h30;
            14'h2624: rddata <= 8'hFB; 14'h2625: rddata <= 8'hC6; 14'h2626: rddata <= 8'h0A; 14'h2627: rddata <= 8'hF5;
            14'h2628: rddata <= 8'h79; 14'h2629: rddata <= 8'hC6; 14'h262A: rddata <= 8'h2F; 14'h262B: rddata <= 8'hCD;
            14'h262C: rddata <= 8'h72; 14'h262D: rddata <= 8'h1D; 14'h262E: rddata <= 8'hF1; 14'h262F: rddata <= 8'hC6;
            14'h2630: rddata <= 8'h30; 14'h2631: rddata <= 8'hCD; 14'h2632: rddata <= 8'h72; 14'h2633: rddata <= 8'h1D;
            14'h2634: rddata <= 8'hC9; 14'h2635: rddata <= 8'h16; 14'h2636: rddata <= 8'h01; 14'h2637: rddata <= 8'h01;
            14'h2638: rddata <= 8'hF0; 14'h2639: rddata <= 8'hD8; 14'h263A: rddata <= 8'hCD; 14'h263B: rddata <= 8'h52;
            14'h263C: rddata <= 8'h26; 14'h263D: rddata <= 8'h01; 14'h263E: rddata <= 8'h18; 14'h263F: rddata <= 8'hFC;
            14'h2640: rddata <= 8'hCD; 14'h2641: rddata <= 8'h52; 14'h2642: rddata <= 8'h26; 14'h2643: rddata <= 8'h01;
            14'h2644: rddata <= 8'h9C; 14'h2645: rddata <= 8'hFF; 14'h2646: rddata <= 8'hCD; 14'h2647: rddata <= 8'h52;
            14'h2648: rddata <= 8'h26; 14'h2649: rddata <= 8'h0E; 14'h264A: rddata <= 8'hF6; 14'h264B: rddata <= 8'hCD;
            14'h264C: rddata <= 8'h52; 14'h264D: rddata <= 8'h26; 14'h264E: rddata <= 8'h16; 14'h264F: rddata <= 8'h00;
            14'h2650: rddata <= 8'h0E; 14'h2651: rddata <= 8'hFF; 14'h2652: rddata <= 8'h3E; 14'h2653: rddata <= 8'hFF;
            14'h2654: rddata <= 8'h3C; 14'h2655: rddata <= 8'h09; 14'h2656: rddata <= 8'h38; 14'h2657: rddata <= 8'hFC;
            14'h2658: rddata <= 8'hED; 14'h2659: rddata <= 8'h42; 14'h265A: rddata <= 8'hB7; 14'h265B: rddata <= 8'h28;
            14'h265C: rddata <= 8'h08; 14'h265D: rddata <= 8'h16; 14'h265E: rddata <= 8'h00; 14'h265F: rddata <= 8'hC6;
            14'h2660: rddata <= 8'h30; 14'h2661: rddata <= 8'hCD; 14'h2662: rddata <= 8'h72; 14'h2663: rddata <= 8'h1D;
            14'h2664: rddata <= 8'hC9; 14'h2665: rddata <= 8'hCB; 14'h2666: rddata <= 8'h42; 14'h2667: rddata <= 8'h28;
            14'h2668: rddata <= 8'hF6; 14'h2669: rddata <= 8'h3E; 14'h266A: rddata <= 8'h20; 14'h266B: rddata <= 8'hCD;
            14'h266C: rddata <= 8'h72; 14'h266D: rddata <= 8'h1D; 14'h266E: rddata <= 8'hC9; 14'h266F: rddata <= 8'h2A;
            14'h2670: rddata <= 8'h4F; 14'h2671: rddata <= 8'h38; 14'h2672: rddata <= 8'h2B; 14'h2673: rddata <= 8'h22;
            14'h2674: rddata <= 8'hCE; 14'h2675: rddata <= 8'h38; 14'h2676: rddata <= 8'h22; 14'h2677: rddata <= 8'hDC;
            14'h2678: rddata <= 8'h38; 14'h2679: rddata <= 8'h2A; 14'h267A: rddata <= 8'hAD; 14'h267B: rddata <= 8'h38;
            14'h267C: rddata <= 8'h22; 14'h267D: rddata <= 8'hC1; 14'h267E: rddata <= 8'h38; 14'h267F: rddata <= 8'h2A;
            14'h2680: rddata <= 8'hD6; 14'h2681: rddata <= 8'h38; 14'h2682: rddata <= 8'h22; 14'h2683: rddata <= 8'hD8;
            14'h2684: rddata <= 8'h38; 14'h2685: rddata <= 8'h22; 14'h2686: rddata <= 8'hDA; 14'h2687: rddata <= 8'h38;
            14'h2688: rddata <= 8'h21; 14'h2689: rddata <= 8'hB1; 14'h268A: rddata <= 8'h38; 14'h268B: rddata <= 8'h22;
            14'h268C: rddata <= 8'hAF; 14'h268D: rddata <= 8'h38; 14'h268E: rddata <= 8'hAF; 14'h268F: rddata <= 8'h6F;
            14'h2690: rddata <= 8'h67; 14'h2691: rddata <= 8'h22; 14'h2692: rddata <= 8'hD4; 14'h2693: rddata <= 8'h38;
            14'h2694: rddata <= 8'h32; 14'h2695: rddata <= 8'hCB; 14'h2696: rddata <= 8'h38; 14'h2697: rddata <= 8'h22;
            14'h2698: rddata <= 8'hDE; 14'h2699: rddata <= 8'h38; 14'h269A: rddata <= 8'hED; 14'h269B: rddata <= 8'h5B;
            14'h269C: rddata <= 8'h4F; 14'h269D: rddata <= 8'h38; 14'h269E: rddata <= 8'h62; 14'h269F: rddata <= 8'h6B;
            14'h26A0: rddata <= 8'h7E; 14'h26A1: rddata <= 8'h23; 14'h26A2: rddata <= 8'hB6; 14'h26A3: rddata <= 8'h28;
            14'h26A4: rddata <= 8'h0E; 14'h26A5: rddata <= 8'h23; 14'h26A6: rddata <= 8'h23; 14'h26A7: rddata <= 8'h23;
            14'h26A8: rddata <= 8'hAF; 14'h26A9: rddata <= 8'hBE; 14'h26AA: rddata <= 8'h23; 14'h26AB: rddata <= 8'h20;
            14'h26AC: rddata <= 8'hFC; 14'h26AD: rddata <= 8'hEB; 14'h26AE: rddata <= 8'h73; 14'h26AF: rddata <= 8'h23;
            14'h26B0: rddata <= 8'h72; 14'h26B1: rddata <= 8'h18; 14'h26B2: rddata <= 8'hEB; 14'h26B3: rddata <= 8'hC9;
            14'h26B4: rddata <= 8'hCD; 14'h26B5: rddata <= 8'h85; 14'h26B6: rddata <= 8'h09; 14'h26B7: rddata <= 8'hE5;
            14'h26B8: rddata <= 8'hCD; 14'h26B9: rddata <= 8'hF7; 14'h26BA: rddata <= 8'h0F; 14'h26BB: rddata <= 8'h32;
            14'h26BC: rddata <= 8'h00; 14'h26BD: rddata <= 8'hBF; 14'h26BE: rddata <= 8'h23; 14'h26BF: rddata <= 8'h23;
            14'h26C0: rddata <= 8'h46; 14'h26C1: rddata <= 8'h23; 14'h26C2: rddata <= 8'h66; 14'h26C3: rddata <= 8'h68;
            14'h26C4: rddata <= 8'h11; 14'h26C5: rddata <= 8'h01; 14'h26C6: rddata <= 8'hBF; 14'h26C7: rddata <= 8'h06;
            14'h26C8: rddata <= 8'h00; 14'h26C9: rddata <= 8'h4F; 14'h26CA: rddata <= 8'hB7; 14'h26CB: rddata <= 8'h28;
            14'h26CC: rddata <= 8'h02; 14'h26CD: rddata <= 8'hED; 14'h26CE: rddata <= 8'hB0; 14'h26CF: rddata <= 8'hAF;
            14'h26D0: rddata <= 8'h12; 14'h26D1: rddata <= 8'hE1; 14'h26D2: rddata <= 8'hC9; 14'h26D3: rddata <= 8'h21;
            14'h26D4: rddata <= 8'h01; 14'h26D5: rddata <= 8'hBF; 14'h26D6: rddata <= 8'h16; 14'h26D7: rddata <= 8'h00;
            14'h26D8: rddata <= 8'h3A; 14'h26D9: rddata <= 8'h00; 14'h26DA: rddata <= 8'hBF; 14'h26DB: rddata <= 8'h3C;
            14'h26DC: rddata <= 8'h5F; 14'h26DD: rddata <= 8'hC3; 14'h26DE: rddata <= 8'h3B; 14'h26DF: rddata <= 8'h27;
            14'h26E0: rddata <= 8'hCD; 14'h26E1: rddata <= 8'h02; 14'h26E2: rddata <= 8'h26; 14'h26E3: rddata <= 8'hB7;
            14'h26E4: rddata <= 8'hFA; 14'h26E5: rddata <= 8'h57; 14'h26E6: rddata <= 8'h25; 14'h26E7: rddata <= 8'hC9;
            14'h26E8: rddata <= 8'h3E; 14'h26E9: rddata <= 8'h1F; 14'h26EA: rddata <= 8'hCD; 14'h26EB: rddata <= 8'hEF;
            14'h26EC: rddata <= 8'h25; 14'h26ED: rddata <= 8'hC3; 14'h26EE: rddata <= 8'hE0; 14'h26EF: rddata <= 8'h26;
            14'h26F0: rddata <= 8'h3E; 14'h26F1: rddata <= 8'h10; 14'h26F2: rddata <= 8'hCD; 14'h26F3: rddata <= 8'hEF;
            14'h26F4: rddata <= 8'h25; 14'h26F5: rddata <= 8'h3E; 14'h26F6: rddata <= 8'h00; 14'h26F7: rddata <= 8'hCD;
            14'h26F8: rddata <= 8'h0B; 14'h26F9: rddata <= 8'h26; 14'h26FA: rddata <= 8'hCD; 14'h26FB: rddata <= 8'hD3;
            14'h26FC: rddata <= 8'h26; 14'h26FD: rddata <= 8'hC3; 14'h26FE: rddata <= 8'hE0; 14'h26FF: rddata <= 8'h26;
            14'h2700: rddata <= 8'h3E; 14'h2701: rddata <= 8'h10; 14'h2702: rddata <= 8'hCD; 14'h2703: rddata <= 8'hEF;
            14'h2704: rddata <= 8'h25; 14'h2705: rddata <= 8'h3E; 14'h2706: rddata <= 8'h19; 14'h2707: rddata <= 8'hCD;
            14'h2708: rddata <= 8'h0B; 14'h2709: rddata <= 8'h26; 14'h270A: rddata <= 8'hCD; 14'h270B: rddata <= 8'hD3;
            14'h270C: rddata <= 8'h26; 14'h270D: rddata <= 8'hC3; 14'h270E: rddata <= 8'hE0; 14'h270F: rddata <= 8'h26;
            14'h2710: rddata <= 8'h3E; 14'h2711: rddata <= 8'h12; 14'h2712: rddata <= 8'hCD; 14'h2713: rddata <= 8'hEF;
            14'h2714: rddata <= 8'h25; 14'h2715: rddata <= 8'hAF; 14'h2716: rddata <= 8'hCD; 14'h2717: rddata <= 8'h0B;
            14'h2718: rddata <= 8'h26; 14'h2719: rddata <= 8'h7B; 14'h271A: rddata <= 8'hCD; 14'h271B: rddata <= 8'h0B;
            14'h271C: rddata <= 8'h26; 14'h271D: rddata <= 8'h7A; 14'h271E: rddata <= 8'hCD; 14'h271F: rddata <= 8'h0B;
            14'h2720: rddata <= 8'h26; 14'h2721: rddata <= 8'hCD; 14'h2722: rddata <= 8'hE0; 14'h2723: rddata <= 8'h26;
            14'h2724: rddata <= 8'hCD; 14'h2725: rddata <= 8'h02; 14'h2726: rddata <= 8'h26; 14'h2727: rddata <= 8'h5F;
            14'h2728: rddata <= 8'hCD; 14'h2729: rddata <= 8'h02; 14'h272A: rddata <= 8'h26; 14'h272B: rddata <= 8'h57;
            14'h272C: rddata <= 8'hD5; 14'h272D: rddata <= 8'h7A; 14'h272E: rddata <= 8'hB3; 14'h272F: rddata <= 8'h28;
            14'h2730: rddata <= 8'h08; 14'h2731: rddata <= 8'hCD; 14'h2732: rddata <= 8'h02; 14'h2733: rddata <= 8'h26;
            14'h2734: rddata <= 8'h77; 14'h2735: rddata <= 8'h23; 14'h2736: rddata <= 8'h1B; 14'h2737: rddata <= 8'h18;
            14'h2738: rddata <= 8'hF4; 14'h2739: rddata <= 8'hD1; 14'h273A: rddata <= 8'hC9; 14'h273B: rddata <= 8'hD5;
            14'h273C: rddata <= 8'h7A; 14'h273D: rddata <= 8'hB3; 14'h273E: rddata <= 8'h28; 14'h273F: rddata <= 8'h08;
            14'h2740: rddata <= 8'h7E; 14'h2741: rddata <= 8'hCD; 14'h2742: rddata <= 8'h0B; 14'h2743: rddata <= 8'h26;
            14'h2744: rddata <= 8'h23; 14'h2745: rddata <= 8'h1B; 14'h2746: rddata <= 8'h18; 14'h2747: rddata <= 8'hF4;
            14'h2748: rddata <= 8'hD1; 14'h2749: rddata <= 8'hC9; 14'h274A: rddata <= 8'h3E; 14'h274B: rddata <= 8'h13;
            14'h274C: rddata <= 8'hCD; 14'h274D: rddata <= 8'hEF; 14'h274E: rddata <= 8'h25; 14'h274F: rddata <= 8'hAF;
            14'h2750: rddata <= 8'hCD; 14'h2751: rddata <= 8'h0B; 14'h2752: rddata <= 8'h26; 14'h2753: rddata <= 8'h7B;
            14'h2754: rddata <= 8'hCD; 14'h2755: rddata <= 8'h0B; 14'h2756: rddata <= 8'h26; 14'h2757: rddata <= 8'h7A;
            14'h2758: rddata <= 8'hCD; 14'h2759: rddata <= 8'h0B; 14'h275A: rddata <= 8'h26; 14'h275B: rddata <= 8'hCD;
            14'h275C: rddata <= 8'h3B; 14'h275D: rddata <= 8'h27; 14'h275E: rddata <= 8'hCD; 14'h275F: rddata <= 8'hE0;
            14'h2760: rddata <= 8'h26; 14'h2761: rddata <= 8'hCD; 14'h2762: rddata <= 8'h02; 14'h2763: rddata <= 8'h26;
            14'h2764: rddata <= 8'h5F; 14'h2765: rddata <= 8'hCD; 14'h2766: rddata <= 8'h02; 14'h2767: rddata <= 8'h26;
            14'h2768: rddata <= 8'h57; 14'h2769: rddata <= 8'hC9; 14'h276A: rddata <= 8'h3E; 14'h276B: rddata <= 8'h14;
            14'h276C: rddata <= 8'hCD; 14'h276D: rddata <= 8'hEF; 14'h276E: rddata <= 8'h25; 14'h276F: rddata <= 8'hAF;
            14'h2770: rddata <= 8'hCD; 14'h2771: rddata <= 8'h0B; 14'h2772: rddata <= 8'h26; 14'h2773: rddata <= 8'h7B;
            14'h2774: rddata <= 8'hCD; 14'h2775: rddata <= 8'h0B; 14'h2776: rddata <= 8'h26; 14'h2777: rddata <= 8'h7A;
            14'h2778: rddata <= 8'hCD; 14'h2779: rddata <= 8'h0B; 14'h277A: rddata <= 8'h26; 14'h277B: rddata <= 8'hAF;
            14'h277C: rddata <= 8'hCD; 14'h277D: rddata <= 8'h0B; 14'h277E: rddata <= 8'h26; 14'h277F: rddata <= 8'hCD;
            14'h2780: rddata <= 8'h0B; 14'h2781: rddata <= 8'h26; 14'h2782: rddata <= 8'hCD; 14'h2783: rddata <= 8'hE0;
            14'h2784: rddata <= 8'h26; 14'h2785: rddata <= 8'hC9; 14'h2786: rddata <= 8'h23; 14'h2787: rddata <= 8'h7E;
            14'h2788: rddata <= 8'hB7; 14'h2789: rddata <= 8'hC8; 14'h278A: rddata <= 8'hFE; 14'h278B: rddata <= 8'h20;
            14'h278C: rddata <= 8'hC0; 14'h278D: rddata <= 8'h18; 14'h278E: rddata <= 8'hF7; 14'h278F: rddata <= 8'h11;
            14'h2790: rddata <= 8'h0D; 14'h2791: rddata <= 8'h00; 14'h2792: rddata <= 8'h21; 14'h2793: rddata <= 8'hEC;
            14'h2794: rddata <= 8'hBF; 14'h2795: rddata <= 8'hCD; 14'h2796: rddata <= 8'h10; 14'h2797: rddata <= 8'h27;
            14'h2798: rddata <= 8'h7B; 14'h2799: rddata <= 8'hFE; 14'h279A: rddata <= 8'h0D; 14'h279B: rddata <= 8'hC2;
            14'h279C: rddata <= 8'hDD; 14'h279D: rddata <= 8'h25; 14'h279E: rddata <= 8'h0E; 14'h279F: rddata <= 8'h0C;
            14'h27A0: rddata <= 8'h21; 14'h27A1: rddata <= 8'hEC; 14'h27A2: rddata <= 8'hBF; 14'h27A3: rddata <= 8'h7E;
            14'h27A4: rddata <= 8'hFE; 14'h27A5: rddata <= 8'hFF; 14'h27A6: rddata <= 8'hC2; 14'h27A7: rddata <= 8'hDD;
            14'h27A8: rddata <= 8'h25; 14'h27A9: rddata <= 8'h23; 14'h27AA: rddata <= 8'h0D; 14'h27AB: rddata <= 8'h20;
            14'h27AC: rddata <= 8'hF6; 14'h27AD: rddata <= 8'h7E; 14'h27AE: rddata <= 8'hB7; 14'h27AF: rddata <= 8'hC2;
            14'h27B0: rddata <= 8'hDD; 14'h27B1: rddata <= 8'h25; 14'h27B2: rddata <= 8'hC9; 14'h27B3: rddata <= 8'hE5;
            14'h27B4: rddata <= 8'hCD; 14'h27B5: rddata <= 8'hF0; 14'h27B6: rddata <= 8'h26; 14'h27B7: rddata <= 8'h2A;
            14'h27B8: rddata <= 8'hFC; 14'h27B9: rddata <= 8'hBF; 14'h27BA: rddata <= 8'h11; 14'h27BB: rddata <= 8'hFF;
            14'h27BC: rddata <= 8'hFF; 14'h27BD: rddata <= 8'hCD; 14'h27BE: rddata <= 8'h10; 14'h27BF: rddata <= 8'h27;
            14'h27C0: rddata <= 8'hCD; 14'h27C1: rddata <= 8'hE8; 14'h27C2: rddata <= 8'h26; 14'h27C3: rddata <= 8'hE1;
            14'h27C4: rddata <= 8'hC9; 14'h27C5: rddata <= 8'hE5; 14'h27C6: rddata <= 8'hCD; 14'h27C7: rddata <= 8'hF0;
            14'h27C8: rddata <= 8'h26; 14'h27C9: rddata <= 8'hCD; 14'h27CA: rddata <= 8'h8F; 14'h27CB: rddata <= 8'h27;
            14'h27CC: rddata <= 8'h11; 14'h27CD: rddata <= 8'h06; 14'h27CE: rddata <= 8'h00; 14'h27CF: rddata <= 8'h21;
            14'h27D0: rddata <= 8'hEC; 14'h27D1: rddata <= 8'hBF; 14'h27D2: rddata <= 8'hCD; 14'h27D3: rddata <= 8'h10;
            14'h27D4: rddata <= 8'h27; 14'h27D5: rddata <= 8'h0E; 14'h27D6: rddata <= 8'h06; 14'h27D7: rddata <= 8'h21;
            14'h27D8: rddata <= 8'hEC; 14'h27D9: rddata <= 8'hBF; 14'h27DA: rddata <= 8'h7E; 14'h27DB: rddata <= 8'hFE;
            14'h27DC: rddata <= 8'h23; 14'h27DD: rddata <= 8'hC2; 14'h27DE: rddata <= 8'hDD; 14'h27DF: rddata <= 8'h25;
            14'h27E0: rddata <= 8'h23; 14'h27E1: rddata <= 8'h0D; 14'h27E2: rddata <= 8'h20; 14'h27E3: rddata <= 8'hF6;
            14'h27E4: rddata <= 8'h2A; 14'h27E5: rddata <= 8'hFC; 14'h27E6: rddata <= 8'hBF; 14'h27E7: rddata <= 8'hED;
            14'h27E8: rddata <= 8'h5B; 14'h27E9: rddata <= 8'hFE; 14'h27EA: rddata <= 8'hBF; 14'h27EB: rddata <= 8'hCD;
            14'h27EC: rddata <= 8'h10; 14'h27ED: rddata <= 8'h27; 14'h27EE: rddata <= 8'hCD; 14'h27EF: rddata <= 8'hE8;
            14'h27F0: rddata <= 8'h26; 14'h27F1: rddata <= 8'hE1; 14'h27F2: rddata <= 8'hC9; 14'h27F3: rddata <= 8'hE5;
            14'h27F4: rddata <= 8'hCD; 14'h27F5: rddata <= 8'hF0; 14'h27F6: rddata <= 8'h26; 14'h27F7: rddata <= 8'hCD;
            14'h27F8: rddata <= 8'h8F; 14'h27F9: rddata <= 8'h27; 14'h27FA: rddata <= 8'h11; 14'h27FB: rddata <= 8'h06;
            14'h27FC: rddata <= 8'h00; 14'h27FD: rddata <= 8'h21; 14'h27FE: rddata <= 8'hEC; 14'h27FF: rddata <= 8'hBF;
            14'h2800: rddata <= 8'hCD; 14'h2801: rddata <= 8'h10; 14'h2802: rddata <= 8'h27; 14'h2803: rddata <= 8'hCD;
            14'h2804: rddata <= 8'h8F; 14'h2805: rddata <= 8'h27; 14'h2806: rddata <= 8'h2A; 14'h2807: rddata <= 8'h4F;
            14'h2808: rddata <= 8'h38; 14'h2809: rddata <= 8'h11; 14'h280A: rddata <= 8'hFF; 14'h280B: rddata <= 8'hFF;
            14'h280C: rddata <= 8'hCD; 14'h280D: rddata <= 8'h10; 14'h280E: rddata <= 8'h27; 14'h280F: rddata <= 8'hCD;
            14'h2810: rddata <= 8'hE8; 14'h2811: rddata <= 8'h26; 14'h2812: rddata <= 8'h2B; 14'h2813: rddata <= 8'hAF;
            14'h2814: rddata <= 8'hBE; 14'h2815: rddata <= 8'h28; 14'h2816: rddata <= 8'hFB; 14'h2817: rddata <= 8'h23;
            14'h2818: rddata <= 8'h23; 14'h2819: rddata <= 8'h23; 14'h281A: rddata <= 8'h23; 14'h281B: rddata <= 8'h22;
            14'h281C: rddata <= 8'hD6; 14'h281D: rddata <= 8'h38; 14'h281E: rddata <= 8'hCD; 14'h281F: rddata <= 8'h6F;
            14'h2820: rddata <= 8'h26; 14'h2821: rddata <= 8'hE1; 14'h2822: rddata <= 8'hC9; 14'h2823: rddata <= 8'hFF;
            14'h2824: rddata <= 8'hFF; 14'h2825: rddata <= 8'hFF; 14'h2826: rddata <= 8'hFF; 14'h2827: rddata <= 8'hFF;
            14'h2828: rddata <= 8'hFF; 14'h2829: rddata <= 8'hFF; 14'h282A: rddata <= 8'hFF; 14'h282B: rddata <= 8'hFF;
            14'h282C: rddata <= 8'hFF; 14'h282D: rddata <= 8'hFF; 14'h282E: rddata <= 8'hFF; 14'h282F: rddata <= 8'h00;
            14'h2830: rddata <= 8'hE5; 14'h2831: rddata <= 8'hCD; 14'h2832: rddata <= 8'h00; 14'h2833: rddata <= 8'h27;
            14'h2834: rddata <= 8'h21; 14'h2835: rddata <= 8'h23; 14'h2836: rddata <= 8'h28; 14'h2837: rddata <= 8'h11;
            14'h2838: rddata <= 8'h0D; 14'h2839: rddata <= 8'h00; 14'h283A: rddata <= 8'hCD; 14'h283B: rddata <= 8'h4A;
            14'h283C: rddata <= 8'h27; 14'h283D: rddata <= 8'h21; 14'h283E: rddata <= 8'h61; 14'h283F: rddata <= 8'h28;
            14'h2840: rddata <= 8'h11; 14'h2841: rddata <= 8'h06; 14'h2842: rddata <= 8'h00; 14'h2843: rddata <= 8'hCD;
            14'h2844: rddata <= 8'h4A; 14'h2845: rddata <= 8'h27; 14'h2846: rddata <= 8'h21; 14'h2847: rddata <= 8'h23;
            14'h2848: rddata <= 8'h28; 14'h2849: rddata <= 8'h11; 14'h284A: rddata <= 8'h0D; 14'h284B: rddata <= 8'h00;
            14'h284C: rddata <= 8'hCD; 14'h284D: rddata <= 8'h4A; 14'h284E: rddata <= 8'h27; 14'h284F: rddata <= 8'hED;
            14'h2850: rddata <= 8'h5B; 14'h2851: rddata <= 8'h4F; 14'h2852: rddata <= 8'h38; 14'h2853: rddata <= 8'h2A;
            14'h2854: rddata <= 8'hD6; 14'h2855: rddata <= 8'h38; 14'h2856: rddata <= 8'hED; 14'h2857: rddata <= 8'h52;
            14'h2858: rddata <= 8'hEB; 14'h2859: rddata <= 8'hCD; 14'h285A: rddata <= 8'h4A; 14'h285B: rddata <= 8'h27;
            14'h285C: rddata <= 8'hCD; 14'h285D: rddata <= 8'hE8; 14'h285E: rddata <= 8'h26; 14'h285F: rddata <= 8'hE1;
            14'h2860: rddata <= 8'hC9; 14'h2861: rddata <= 8'h42; 14'h2862: rddata <= 8'h41; 14'h2863: rddata <= 8'h53;
            14'h2864: rddata <= 8'h50; 14'h2865: rddata <= 8'h52; 14'h2866: rddata <= 8'h47; 14'h2867: rddata <= 8'hE5;
            14'h2868: rddata <= 8'hCD; 14'h2869: rddata <= 8'h00; 14'h286A: rddata <= 8'h27; 14'h286B: rddata <= 8'h21;
            14'h286C: rddata <= 8'h23; 14'h286D: rddata <= 8'h28; 14'h286E: rddata <= 8'h11; 14'h286F: rddata <= 8'h0D;
            14'h2870: rddata <= 8'h00; 14'h2871: rddata <= 8'hCD; 14'h2872: rddata <= 8'h4A; 14'h2873: rddata <= 8'h27;
            14'h2874: rddata <= 8'h21; 14'h2875: rddata <= 8'h8C; 14'h2876: rddata <= 8'h28; 14'h2877: rddata <= 8'h11;
            14'h2878: rddata <= 8'h06; 14'h2879: rddata <= 8'h00; 14'h287A: rddata <= 8'hCD; 14'h287B: rddata <= 8'h4A;
            14'h287C: rddata <= 8'h27; 14'h287D: rddata <= 8'h2A; 14'h287E: rddata <= 8'hFC; 14'h287F: rddata <= 8'hBF;
            14'h2880: rddata <= 8'hED; 14'h2881: rddata <= 8'h5B; 14'h2882: rddata <= 8'hFE; 14'h2883: rddata <= 8'hBF;
            14'h2884: rddata <= 8'hCD; 14'h2885: rddata <= 8'h4A; 14'h2886: rddata <= 8'h27; 14'h2887: rddata <= 8'hCD;
            14'h2888: rddata <= 8'hE8; 14'h2889: rddata <= 8'h26; 14'h288A: rddata <= 8'hE1; 14'h288B: rddata <= 8'hC9;
            14'h288C: rddata <= 8'h23; 14'h288D: rddata <= 8'h23; 14'h288E: rddata <= 8'h23; 14'h288F: rddata <= 8'h23;
            14'h2890: rddata <= 8'h23; 14'h2891: rddata <= 8'h23; 14'h2892: rddata <= 8'hE5; 14'h2893: rddata <= 8'hCD;
            14'h2894: rddata <= 8'h00; 14'h2895: rddata <= 8'h27; 14'h2896: rddata <= 8'h2A; 14'h2897: rddata <= 8'hFC;
            14'h2898: rddata <= 8'hBF; 14'h2899: rddata <= 8'hED; 14'h289A: rddata <= 8'h5B; 14'h289B: rddata <= 8'hFE;
            14'h289C: rddata <= 8'hBF; 14'h289D: rddata <= 8'hCD; 14'h289E: rddata <= 8'h4A; 14'h289F: rddata <= 8'h27;
            14'h28A0: rddata <= 8'hCD; 14'h28A1: rddata <= 8'hE8; 14'h28A2: rddata <= 8'h26; 14'h28A3: rddata <= 8'hE1;
            14'h28A4: rddata <= 8'hC9; 14'h28A5: rddata <= 8'hCD; 14'h28A6: rddata <= 8'hE8; 14'h28A7: rddata <= 8'h26;
            14'h28A8: rddata <= 8'hCD; 14'h28A9: rddata <= 8'hB4; 14'h28AA: rddata <= 8'h26; 14'h28AB: rddata <= 8'h3A;
            14'h28AC: rddata <= 8'h00; 14'h28AD: rddata <= 8'hBF; 14'h28AE: rddata <= 8'hFE; 14'h28AF: rddata <= 8'h05;
            14'h28B0: rddata <= 8'h38; 14'h28B1: rddata <= 8'h0D; 14'h28B2: rddata <= 8'hD6; 14'h28B3: rddata <= 8'h03;
            14'h28B4: rddata <= 8'h16; 14'h28B5: rddata <= 8'hBF; 14'h28B6: rddata <= 8'h5F; 14'h28B7: rddata <= 8'h21;
            14'h28B8: rddata <= 8'hD1; 14'h28B9: rddata <= 8'h28; 14'h28BA: rddata <= 8'hCD; 14'h28BB: rddata <= 8'hC5;
            14'h28BC: rddata <= 8'h28; 14'h28BD: rddata <= 8'h28; 14'h28BE: rddata <= 8'h17; 14'h28BF: rddata <= 8'hCD;
            14'h28C0: rddata <= 8'hF3; 14'h28C1: rddata <= 8'h27; 14'h28C2: rddata <= 8'hC3; 14'h28C3: rddata <= 8'hCB;
            14'h28C4: rddata <= 8'h0B; 14'h28C5: rddata <= 8'h1A; 14'h28C6: rddata <= 8'hCD; 14'h28C7: rddata <= 8'h28;
            14'h28C8: rddata <= 8'h29; 14'h28C9: rddata <= 8'h13; 14'h28CA: rddata <= 8'hBE; 14'h28CB: rddata <= 8'h23;
            14'h28CC: rddata <= 8'hC0; 14'h28CD: rddata <= 8'hB7; 14'h28CE: rddata <= 8'h20; 14'h28CF: rddata <= 8'hF5;
            14'h28D0: rddata <= 8'hC9; 14'h28D1: rddata <= 8'h2E; 14'h28D2: rddata <= 8'h52; 14'h28D3: rddata <= 8'h4F;
            14'h28D4: rddata <= 8'h4D; 14'h28D5: rddata <= 8'h00; 14'h28D6: rddata <= 8'hCD; 14'h28D7: rddata <= 8'hF0;
            14'h28D8: rddata <= 8'h26; 14'h28D9: rddata <= 8'h3E; 14'h28DA: rddata <= 8'h23; 14'h28DB: rddata <= 8'hD3;
            14'h28DC: rddata <= 8'hF3; 14'h28DD: rddata <= 8'h21; 14'h28DE: rddata <= 8'h00; 14'h28DF: rddata <= 8'hC0;
            14'h28E0: rddata <= 8'h11; 14'h28E1: rddata <= 8'h00; 14'h28E2: rddata <= 8'h40; 14'h28E3: rddata <= 8'hCD;
            14'h28E4: rddata <= 8'h10; 14'h28E5: rddata <= 8'h27; 14'h28E6: rddata <= 8'h7A; 14'h28E7: rddata <= 8'hFE;
            14'h28E8: rddata <= 8'h20; 14'h28E9: rddata <= 8'h20; 14'h28EA: rddata <= 8'h0B; 14'h28EB: rddata <= 8'h21;
            14'h28EC: rddata <= 8'h00; 14'h28ED: rddata <= 8'hC0; 14'h28EE: rddata <= 8'h11; 14'h28EF: rddata <= 8'h00;
            14'h28F0: rddata <= 8'hE0; 14'h28F1: rddata <= 8'h01; 14'h28F2: rddata <= 8'h00; 14'h28F3: rddata <= 8'h20;
            14'h28F4: rddata <= 8'hED; 14'h28F5: rddata <= 8'hB0; 14'h28F6: rddata <= 8'hCD; 14'h28F7: rddata <= 8'hE8;
            14'h28F8: rddata <= 8'h26; 14'h28F9: rddata <= 8'hAF; 14'h28FA: rddata <= 8'h21; 14'h28FB: rddata <= 8'h03;
            14'h28FC: rddata <= 8'hE0; 14'h28FD: rddata <= 8'h06; 14'h28FE: rddata <= 8'h0C; 14'h28FF: rddata <= 8'h86;
            14'h2900: rddata <= 8'h23; 14'h2901: rddata <= 8'h80; 14'h2902: rddata <= 8'h05; 14'h2903: rddata <= 8'h20;
            14'h2904: rddata <= 8'hFA; 14'h2905: rddata <= 8'hAE; 14'h2906: rddata <= 8'h47; 14'h2907: rddata <= 8'h21;
            14'h2908: rddata <= 8'h00; 14'h2909: rddata <= 8'hC0; 14'h290A: rddata <= 8'h11; 14'h290B: rddata <= 8'h00;
            14'h290C: rddata <= 8'h40; 14'h290D: rddata <= 8'h78; 14'h290E: rddata <= 8'hAE; 14'h290F: rddata <= 8'h77;
            14'h2910: rddata <= 8'h23; 14'h2911: rddata <= 8'h1B; 14'h2912: rddata <= 8'h7A; 14'h2913: rddata <= 8'hB3;
            14'h2914: rddata <= 8'h20; 14'h2915: rddata <= 8'hF7; 14'h2916: rddata <= 8'h3E; 14'h2917: rddata <= 8'h21;
            14'h2918: rddata <= 8'hD3; 14'h2919: rddata <= 8'hF1; 14'h291A: rddata <= 8'h3E; 14'h291B: rddata <= 8'h22;
            14'h291C: rddata <= 8'hD3; 14'h291D: rddata <= 8'hF2; 14'h291E: rddata <= 8'h3E; 14'h291F: rddata <= 8'hA3;
            14'h2920: rddata <= 8'hD3; 14'h2921: rddata <= 8'hF3; 14'h2922: rddata <= 8'h31; 14'h2923: rddata <= 8'hA0;
            14'h2924: rddata <= 8'h38; 14'h2925: rddata <= 8'hC3; 14'h2926: rddata <= 8'h10; 14'h2927: rddata <= 8'hE0;
            14'h2928: rddata <= 8'hFE; 14'h2929: rddata <= 8'h61; 14'h292A: rddata <= 8'hD8; 14'h292B: rddata <= 8'hFE;
            14'h292C: rddata <= 8'h7B; 14'h292D: rddata <= 8'hD0; 14'h292E: rddata <= 8'hD6; 14'h292F: rddata <= 8'h20;
            14'h2930: rddata <= 8'hC9; 14'h2931: rddata <= 8'hFF; 14'h2932: rddata <= 8'hFF; 14'h2933: rddata <= 8'hFF;
            14'h2934: rddata <= 8'hFF; 14'h2935: rddata <= 8'hFF; 14'h2936: rddata <= 8'hFF; 14'h2937: rddata <= 8'hFF;
            14'h2938: rddata <= 8'hFF; 14'h2939: rddata <= 8'hFF; 14'h293A: rddata <= 8'hFF; 14'h293B: rddata <= 8'hFF;
            14'h293C: rddata <= 8'hFF; 14'h293D: rddata <= 8'hFF; 14'h293E: rddata <= 8'hFF; 14'h293F: rddata <= 8'hFF;
            14'h2940: rddata <= 8'hFF; 14'h2941: rddata <= 8'hFF; 14'h2942: rddata <= 8'hFF; 14'h2943: rddata <= 8'hFF;
            14'h2944: rddata <= 8'hFF; 14'h2945: rddata <= 8'hFF; 14'h2946: rddata <= 8'hFF; 14'h2947: rddata <= 8'hFF;
            14'h2948: rddata <= 8'hFF; 14'h2949: rddata <= 8'hFF; 14'h294A: rddata <= 8'hFF; 14'h294B: rddata <= 8'hFF;
            14'h294C: rddata <= 8'hFF; 14'h294D: rddata <= 8'hFF; 14'h294E: rddata <= 8'hFF; 14'h294F: rddata <= 8'hFF;
            14'h2950: rddata <= 8'hFF; 14'h2951: rddata <= 8'hFF; 14'h2952: rddata <= 8'hFF; 14'h2953: rddata <= 8'hFF;
            14'h2954: rddata <= 8'hFF; 14'h2955: rddata <= 8'hFF; 14'h2956: rddata <= 8'hFF; 14'h2957: rddata <= 8'hFF;
            14'h2958: rddata <= 8'hFF; 14'h2959: rddata <= 8'hFF; 14'h295A: rddata <= 8'hFF; 14'h295B: rddata <= 8'hFF;
            14'h295C: rddata <= 8'hFF; 14'h295D: rddata <= 8'hFF; 14'h295E: rddata <= 8'hFF; 14'h295F: rddata <= 8'hFF;
            14'h2960: rddata <= 8'hFF; 14'h2961: rddata <= 8'hFF; 14'h2962: rddata <= 8'hFF; 14'h2963: rddata <= 8'hFF;
            14'h2964: rddata <= 8'hFF; 14'h2965: rddata <= 8'hFF; 14'h2966: rddata <= 8'hFF; 14'h2967: rddata <= 8'hFF;
            14'h2968: rddata <= 8'hFF; 14'h2969: rddata <= 8'hFF; 14'h296A: rddata <= 8'hFF; 14'h296B: rddata <= 8'hFF;
            14'h296C: rddata <= 8'hFF; 14'h296D: rddata <= 8'hFF; 14'h296E: rddata <= 8'hFF; 14'h296F: rddata <= 8'hFF;
            14'h2970: rddata <= 8'hFF; 14'h2971: rddata <= 8'hFF; 14'h2972: rddata <= 8'hFF; 14'h2973: rddata <= 8'hFF;
            14'h2974: rddata <= 8'hFF; 14'h2975: rddata <= 8'hFF; 14'h2976: rddata <= 8'hFF; 14'h2977: rddata <= 8'hFF;
            14'h2978: rddata <= 8'hFF; 14'h2979: rddata <= 8'hFF; 14'h297A: rddata <= 8'hFF; 14'h297B: rddata <= 8'hFF;
            14'h297C: rddata <= 8'hFF; 14'h297D: rddata <= 8'hFF; 14'h297E: rddata <= 8'hFF; 14'h297F: rddata <= 8'hFF;
            14'h2980: rddata <= 8'hFF; 14'h2981: rddata <= 8'hFF; 14'h2982: rddata <= 8'hFF; 14'h2983: rddata <= 8'hFF;
            14'h2984: rddata <= 8'hFF; 14'h2985: rddata <= 8'hFF; 14'h2986: rddata <= 8'hFF; 14'h2987: rddata <= 8'hFF;
            14'h2988: rddata <= 8'hFF; 14'h2989: rddata <= 8'hFF; 14'h298A: rddata <= 8'hFF; 14'h298B: rddata <= 8'hFF;
            14'h298C: rddata <= 8'hFF; 14'h298D: rddata <= 8'hFF; 14'h298E: rddata <= 8'hFF; 14'h298F: rddata <= 8'hFF;
            14'h2990: rddata <= 8'hFF; 14'h2991: rddata <= 8'hFF; 14'h2992: rddata <= 8'hFF; 14'h2993: rddata <= 8'hFF;
            14'h2994: rddata <= 8'hFF; 14'h2995: rddata <= 8'hFF; 14'h2996: rddata <= 8'hFF; 14'h2997: rddata <= 8'hFF;
            14'h2998: rddata <= 8'hFF; 14'h2999: rddata <= 8'hFF; 14'h299A: rddata <= 8'hFF; 14'h299B: rddata <= 8'hFF;
            14'h299C: rddata <= 8'hFF; 14'h299D: rddata <= 8'hFF; 14'h299E: rddata <= 8'hFF; 14'h299F: rddata <= 8'hFF;
            14'h29A0: rddata <= 8'hFF; 14'h29A1: rddata <= 8'hFF; 14'h29A2: rddata <= 8'hFF; 14'h29A3: rddata <= 8'hFF;
            14'h29A4: rddata <= 8'hFF; 14'h29A5: rddata <= 8'hFF; 14'h29A6: rddata <= 8'hFF; 14'h29A7: rddata <= 8'hFF;
            14'h29A8: rddata <= 8'hFF; 14'h29A9: rddata <= 8'hFF; 14'h29AA: rddata <= 8'hFF; 14'h29AB: rddata <= 8'hFF;
            14'h29AC: rddata <= 8'hFF; 14'h29AD: rddata <= 8'hFF; 14'h29AE: rddata <= 8'hFF; 14'h29AF: rddata <= 8'hFF;
            14'h29B0: rddata <= 8'hFF; 14'h29B1: rddata <= 8'hFF; 14'h29B2: rddata <= 8'hFF; 14'h29B3: rddata <= 8'hFF;
            14'h29B4: rddata <= 8'hFF; 14'h29B5: rddata <= 8'hFF; 14'h29B6: rddata <= 8'hFF; 14'h29B7: rddata <= 8'hFF;
            14'h29B8: rddata <= 8'hFF; 14'h29B9: rddata <= 8'hFF; 14'h29BA: rddata <= 8'hFF; 14'h29BB: rddata <= 8'hFF;
            14'h29BC: rddata <= 8'hFF; 14'h29BD: rddata <= 8'hFF; 14'h29BE: rddata <= 8'hFF; 14'h29BF: rddata <= 8'hFF;
            14'h29C0: rddata <= 8'hFF; 14'h29C1: rddata <= 8'hFF; 14'h29C2: rddata <= 8'hFF; 14'h29C3: rddata <= 8'hFF;
            14'h29C4: rddata <= 8'hFF; 14'h29C5: rddata <= 8'hFF; 14'h29C6: rddata <= 8'hFF; 14'h29C7: rddata <= 8'hFF;
            14'h29C8: rddata <= 8'hFF; 14'h29C9: rddata <= 8'hFF; 14'h29CA: rddata <= 8'hFF; 14'h29CB: rddata <= 8'hFF;
            14'h29CC: rddata <= 8'hFF; 14'h29CD: rddata <= 8'hFF; 14'h29CE: rddata <= 8'hFF; 14'h29CF: rddata <= 8'hFF;
            14'h29D0: rddata <= 8'hFF; 14'h29D1: rddata <= 8'hFF; 14'h29D2: rddata <= 8'hFF; 14'h29D3: rddata <= 8'hFF;
            14'h29D4: rddata <= 8'hFF; 14'h29D5: rddata <= 8'hFF; 14'h29D6: rddata <= 8'hFF; 14'h29D7: rddata <= 8'hFF;
            14'h29D8: rddata <= 8'hFF; 14'h29D9: rddata <= 8'hFF; 14'h29DA: rddata <= 8'hFF; 14'h29DB: rddata <= 8'hFF;
            14'h29DC: rddata <= 8'hFF; 14'h29DD: rddata <= 8'hFF; 14'h29DE: rddata <= 8'hFF; 14'h29DF: rddata <= 8'hFF;
            14'h29E0: rddata <= 8'hFF; 14'h29E1: rddata <= 8'hFF; 14'h29E2: rddata <= 8'hFF; 14'h29E3: rddata <= 8'hFF;
            14'h29E4: rddata <= 8'hFF; 14'h29E5: rddata <= 8'hFF; 14'h29E6: rddata <= 8'hFF; 14'h29E7: rddata <= 8'hFF;
            14'h29E8: rddata <= 8'hFF; 14'h29E9: rddata <= 8'hFF; 14'h29EA: rddata <= 8'hFF; 14'h29EB: rddata <= 8'hFF;
            14'h29EC: rddata <= 8'hFF; 14'h29ED: rddata <= 8'hFF; 14'h29EE: rddata <= 8'hFF; 14'h29EF: rddata <= 8'hFF;
            14'h29F0: rddata <= 8'hFF; 14'h29F1: rddata <= 8'hFF; 14'h29F2: rddata <= 8'hFF; 14'h29F3: rddata <= 8'hFF;
            14'h29F4: rddata <= 8'hFF; 14'h29F5: rddata <= 8'hFF; 14'h29F6: rddata <= 8'hFF; 14'h29F7: rddata <= 8'hFF;
            14'h29F8: rddata <= 8'hFF; 14'h29F9: rddata <= 8'hFF; 14'h29FA: rddata <= 8'hFF; 14'h29FB: rddata <= 8'hFF;
            14'h29FC: rddata <= 8'hFF; 14'h29FD: rddata <= 8'hFF; 14'h29FE: rddata <= 8'hFF; 14'h29FF: rddata <= 8'hFF;
            14'h2A00: rddata <= 8'hFF; 14'h2A01: rddata <= 8'hFF; 14'h2A02: rddata <= 8'hFF; 14'h2A03: rddata <= 8'hFF;
            14'h2A04: rddata <= 8'hFF; 14'h2A05: rddata <= 8'hFF; 14'h2A06: rddata <= 8'hFF; 14'h2A07: rddata <= 8'hFF;
            14'h2A08: rddata <= 8'hFF; 14'h2A09: rddata <= 8'hFF; 14'h2A0A: rddata <= 8'hFF; 14'h2A0B: rddata <= 8'hFF;
            14'h2A0C: rddata <= 8'hFF; 14'h2A0D: rddata <= 8'hFF; 14'h2A0E: rddata <= 8'hFF; 14'h2A0F: rddata <= 8'hFF;
            14'h2A10: rddata <= 8'hFF; 14'h2A11: rddata <= 8'hFF; 14'h2A12: rddata <= 8'hFF; 14'h2A13: rddata <= 8'hFF;
            14'h2A14: rddata <= 8'hFF; 14'h2A15: rddata <= 8'hFF; 14'h2A16: rddata <= 8'hFF; 14'h2A17: rddata <= 8'hFF;
            14'h2A18: rddata <= 8'hFF; 14'h2A19: rddata <= 8'hFF; 14'h2A1A: rddata <= 8'hFF; 14'h2A1B: rddata <= 8'hFF;
            14'h2A1C: rddata <= 8'hFF; 14'h2A1D: rddata <= 8'hFF; 14'h2A1E: rddata <= 8'hFF; 14'h2A1F: rddata <= 8'hFF;
            14'h2A20: rddata <= 8'hFF; 14'h2A21: rddata <= 8'hFF; 14'h2A22: rddata <= 8'hFF; 14'h2A23: rddata <= 8'hFF;
            14'h2A24: rddata <= 8'hFF; 14'h2A25: rddata <= 8'hFF; 14'h2A26: rddata <= 8'hFF; 14'h2A27: rddata <= 8'hFF;
            14'h2A28: rddata <= 8'hFF; 14'h2A29: rddata <= 8'hFF; 14'h2A2A: rddata <= 8'hFF; 14'h2A2B: rddata <= 8'hFF;
            14'h2A2C: rddata <= 8'hFF; 14'h2A2D: rddata <= 8'hFF; 14'h2A2E: rddata <= 8'hFF; 14'h2A2F: rddata <= 8'hFF;
            14'h2A30: rddata <= 8'hFF; 14'h2A31: rddata <= 8'hFF; 14'h2A32: rddata <= 8'hFF; 14'h2A33: rddata <= 8'hFF;
            14'h2A34: rddata <= 8'hFF; 14'h2A35: rddata <= 8'hFF; 14'h2A36: rddata <= 8'hFF; 14'h2A37: rddata <= 8'hFF;
            14'h2A38: rddata <= 8'hFF; 14'h2A39: rddata <= 8'hFF; 14'h2A3A: rddata <= 8'hFF; 14'h2A3B: rddata <= 8'hFF;
            14'h2A3C: rddata <= 8'hFF; 14'h2A3D: rddata <= 8'hFF; 14'h2A3E: rddata <= 8'hFF; 14'h2A3F: rddata <= 8'hFF;
            14'h2A40: rddata <= 8'hFF; 14'h2A41: rddata <= 8'hFF; 14'h2A42: rddata <= 8'hFF; 14'h2A43: rddata <= 8'hFF;
            14'h2A44: rddata <= 8'hFF; 14'h2A45: rddata <= 8'hFF; 14'h2A46: rddata <= 8'hFF; 14'h2A47: rddata <= 8'hFF;
            14'h2A48: rddata <= 8'hFF; 14'h2A49: rddata <= 8'hFF; 14'h2A4A: rddata <= 8'hFF; 14'h2A4B: rddata <= 8'hFF;
            14'h2A4C: rddata <= 8'hFF; 14'h2A4D: rddata <= 8'hFF; 14'h2A4E: rddata <= 8'hFF; 14'h2A4F: rddata <= 8'hFF;
            14'h2A50: rddata <= 8'hFF; 14'h2A51: rddata <= 8'hFF; 14'h2A52: rddata <= 8'hFF; 14'h2A53: rddata <= 8'hFF;
            14'h2A54: rddata <= 8'hFF; 14'h2A55: rddata <= 8'hFF; 14'h2A56: rddata <= 8'hFF; 14'h2A57: rddata <= 8'hFF;
            14'h2A58: rddata <= 8'hFF; 14'h2A59: rddata <= 8'hFF; 14'h2A5A: rddata <= 8'hFF; 14'h2A5B: rddata <= 8'hFF;
            14'h2A5C: rddata <= 8'hFF; 14'h2A5D: rddata <= 8'hFF; 14'h2A5E: rddata <= 8'hFF; 14'h2A5F: rddata <= 8'hFF;
            14'h2A60: rddata <= 8'hFF; 14'h2A61: rddata <= 8'hFF; 14'h2A62: rddata <= 8'hFF; 14'h2A63: rddata <= 8'hFF;
            14'h2A64: rddata <= 8'hFF; 14'h2A65: rddata <= 8'hFF; 14'h2A66: rddata <= 8'hFF; 14'h2A67: rddata <= 8'hFF;
            14'h2A68: rddata <= 8'hFF; 14'h2A69: rddata <= 8'hFF; 14'h2A6A: rddata <= 8'hFF; 14'h2A6B: rddata <= 8'hFF;
            14'h2A6C: rddata <= 8'hFF; 14'h2A6D: rddata <= 8'hFF; 14'h2A6E: rddata <= 8'hFF; 14'h2A6F: rddata <= 8'hFF;
            14'h2A70: rddata <= 8'hFF; 14'h2A71: rddata <= 8'hFF; 14'h2A72: rddata <= 8'hFF; 14'h2A73: rddata <= 8'hFF;
            14'h2A74: rddata <= 8'hFF; 14'h2A75: rddata <= 8'hFF; 14'h2A76: rddata <= 8'hFF; 14'h2A77: rddata <= 8'hFF;
            14'h2A78: rddata <= 8'hFF; 14'h2A79: rddata <= 8'hFF; 14'h2A7A: rddata <= 8'hFF; 14'h2A7B: rddata <= 8'hFF;
            14'h2A7C: rddata <= 8'hFF; 14'h2A7D: rddata <= 8'hFF; 14'h2A7E: rddata <= 8'hFF; 14'h2A7F: rddata <= 8'hFF;
            14'h2A80: rddata <= 8'hFF; 14'h2A81: rddata <= 8'hFF; 14'h2A82: rddata <= 8'hFF; 14'h2A83: rddata <= 8'hFF;
            14'h2A84: rddata <= 8'hFF; 14'h2A85: rddata <= 8'hFF; 14'h2A86: rddata <= 8'hFF; 14'h2A87: rddata <= 8'hFF;
            14'h2A88: rddata <= 8'hFF; 14'h2A89: rddata <= 8'hFF; 14'h2A8A: rddata <= 8'hFF; 14'h2A8B: rddata <= 8'hFF;
            14'h2A8C: rddata <= 8'hFF; 14'h2A8D: rddata <= 8'hFF; 14'h2A8E: rddata <= 8'hFF; 14'h2A8F: rddata <= 8'hFF;
            14'h2A90: rddata <= 8'hFF; 14'h2A91: rddata <= 8'hFF; 14'h2A92: rddata <= 8'hFF; 14'h2A93: rddata <= 8'hFF;
            14'h2A94: rddata <= 8'hFF; 14'h2A95: rddata <= 8'hFF; 14'h2A96: rddata <= 8'hFF; 14'h2A97: rddata <= 8'hFF;
            14'h2A98: rddata <= 8'hFF; 14'h2A99: rddata <= 8'hFF; 14'h2A9A: rddata <= 8'hFF; 14'h2A9B: rddata <= 8'hFF;
            14'h2A9C: rddata <= 8'hFF; 14'h2A9D: rddata <= 8'hFF; 14'h2A9E: rddata <= 8'hFF; 14'h2A9F: rddata <= 8'hFF;
            14'h2AA0: rddata <= 8'hFF; 14'h2AA1: rddata <= 8'hFF; 14'h2AA2: rddata <= 8'hFF; 14'h2AA3: rddata <= 8'hFF;
            14'h2AA4: rddata <= 8'hFF; 14'h2AA5: rddata <= 8'hFF; 14'h2AA6: rddata <= 8'hFF; 14'h2AA7: rddata <= 8'hFF;
            14'h2AA8: rddata <= 8'hFF; 14'h2AA9: rddata <= 8'hFF; 14'h2AAA: rddata <= 8'hFF; 14'h2AAB: rddata <= 8'hFF;
            14'h2AAC: rddata <= 8'hFF; 14'h2AAD: rddata <= 8'hFF; 14'h2AAE: rddata <= 8'hFF; 14'h2AAF: rddata <= 8'hFF;
            14'h2AB0: rddata <= 8'hFF; 14'h2AB1: rddata <= 8'hFF; 14'h2AB2: rddata <= 8'hFF; 14'h2AB3: rddata <= 8'hFF;
            14'h2AB4: rddata <= 8'hFF; 14'h2AB5: rddata <= 8'hFF; 14'h2AB6: rddata <= 8'hFF; 14'h2AB7: rddata <= 8'hFF;
            14'h2AB8: rddata <= 8'hFF; 14'h2AB9: rddata <= 8'hFF; 14'h2ABA: rddata <= 8'hFF; 14'h2ABB: rddata <= 8'hFF;
            14'h2ABC: rddata <= 8'hFF; 14'h2ABD: rddata <= 8'hFF; 14'h2ABE: rddata <= 8'hFF; 14'h2ABF: rddata <= 8'hFF;
            14'h2AC0: rddata <= 8'hFF; 14'h2AC1: rddata <= 8'hFF; 14'h2AC2: rddata <= 8'hFF; 14'h2AC3: rddata <= 8'hFF;
            14'h2AC4: rddata <= 8'hFF; 14'h2AC5: rddata <= 8'hFF; 14'h2AC6: rddata <= 8'hFF; 14'h2AC7: rddata <= 8'hFF;
            14'h2AC8: rddata <= 8'hFF; 14'h2AC9: rddata <= 8'hFF; 14'h2ACA: rddata <= 8'hFF; 14'h2ACB: rddata <= 8'hFF;
            14'h2ACC: rddata <= 8'hFF; 14'h2ACD: rddata <= 8'hFF; 14'h2ACE: rddata <= 8'hFF; 14'h2ACF: rddata <= 8'hFF;
            14'h2AD0: rddata <= 8'hFF; 14'h2AD1: rddata <= 8'hFF; 14'h2AD2: rddata <= 8'hFF; 14'h2AD3: rddata <= 8'hFF;
            14'h2AD4: rddata <= 8'hFF; 14'h2AD5: rddata <= 8'hFF; 14'h2AD6: rddata <= 8'hFF; 14'h2AD7: rddata <= 8'hFF;
            14'h2AD8: rddata <= 8'hFF; 14'h2AD9: rddata <= 8'hFF; 14'h2ADA: rddata <= 8'hFF; 14'h2ADB: rddata <= 8'hFF;
            14'h2ADC: rddata <= 8'hFF; 14'h2ADD: rddata <= 8'hFF; 14'h2ADE: rddata <= 8'hFF; 14'h2ADF: rddata <= 8'hFF;
            14'h2AE0: rddata <= 8'hFF; 14'h2AE1: rddata <= 8'hFF; 14'h2AE2: rddata <= 8'hFF; 14'h2AE3: rddata <= 8'hFF;
            14'h2AE4: rddata <= 8'hFF; 14'h2AE5: rddata <= 8'hFF; 14'h2AE6: rddata <= 8'hFF; 14'h2AE7: rddata <= 8'hFF;
            14'h2AE8: rddata <= 8'hFF; 14'h2AE9: rddata <= 8'hFF; 14'h2AEA: rddata <= 8'hFF; 14'h2AEB: rddata <= 8'hFF;
            14'h2AEC: rddata <= 8'hFF; 14'h2AED: rddata <= 8'hFF; 14'h2AEE: rddata <= 8'hFF; 14'h2AEF: rddata <= 8'hFF;
            14'h2AF0: rddata <= 8'hFF; 14'h2AF1: rddata <= 8'hFF; 14'h2AF2: rddata <= 8'hFF; 14'h2AF3: rddata <= 8'hFF;
            14'h2AF4: rddata <= 8'hFF; 14'h2AF5: rddata <= 8'hFF; 14'h2AF6: rddata <= 8'hFF; 14'h2AF7: rddata <= 8'hFF;
            14'h2AF8: rddata <= 8'hFF; 14'h2AF9: rddata <= 8'hFF; 14'h2AFA: rddata <= 8'hFF; 14'h2AFB: rddata <= 8'hFF;
            14'h2AFC: rddata <= 8'hFF; 14'h2AFD: rddata <= 8'hFF; 14'h2AFE: rddata <= 8'hFF; 14'h2AFF: rddata <= 8'hFF;
            14'h2B00: rddata <= 8'hFF; 14'h2B01: rddata <= 8'hFF; 14'h2B02: rddata <= 8'hFF; 14'h2B03: rddata <= 8'hFF;
            14'h2B04: rddata <= 8'hFF; 14'h2B05: rddata <= 8'hFF; 14'h2B06: rddata <= 8'hFF; 14'h2B07: rddata <= 8'hFF;
            14'h2B08: rddata <= 8'hFF; 14'h2B09: rddata <= 8'hFF; 14'h2B0A: rddata <= 8'hFF; 14'h2B0B: rddata <= 8'hFF;
            14'h2B0C: rddata <= 8'hFF; 14'h2B0D: rddata <= 8'hFF; 14'h2B0E: rddata <= 8'hFF; 14'h2B0F: rddata <= 8'hFF;
            14'h2B10: rddata <= 8'hFF; 14'h2B11: rddata <= 8'hFF; 14'h2B12: rddata <= 8'hFF; 14'h2B13: rddata <= 8'hFF;
            14'h2B14: rddata <= 8'hFF; 14'h2B15: rddata <= 8'hFF; 14'h2B16: rddata <= 8'hFF; 14'h2B17: rddata <= 8'hFF;
            14'h2B18: rddata <= 8'hFF; 14'h2B19: rddata <= 8'hFF; 14'h2B1A: rddata <= 8'hFF; 14'h2B1B: rddata <= 8'hFF;
            14'h2B1C: rddata <= 8'hFF; 14'h2B1D: rddata <= 8'hFF; 14'h2B1E: rddata <= 8'hFF; 14'h2B1F: rddata <= 8'hFF;
            14'h2B20: rddata <= 8'hFF; 14'h2B21: rddata <= 8'hFF; 14'h2B22: rddata <= 8'hFF; 14'h2B23: rddata <= 8'hFF;
            14'h2B24: rddata <= 8'hFF; 14'h2B25: rddata <= 8'hFF; 14'h2B26: rddata <= 8'hFF; 14'h2B27: rddata <= 8'hFF;
            14'h2B28: rddata <= 8'hFF; 14'h2B29: rddata <= 8'hFF; 14'h2B2A: rddata <= 8'hFF; 14'h2B2B: rddata <= 8'hFF;
            14'h2B2C: rddata <= 8'hFF; 14'h2B2D: rddata <= 8'hFF; 14'h2B2E: rddata <= 8'hFF; 14'h2B2F: rddata <= 8'hFF;
            14'h2B30: rddata <= 8'hFF; 14'h2B31: rddata <= 8'hFF; 14'h2B32: rddata <= 8'hFF; 14'h2B33: rddata <= 8'hFF;
            14'h2B34: rddata <= 8'hFF; 14'h2B35: rddata <= 8'hFF; 14'h2B36: rddata <= 8'hFF; 14'h2B37: rddata <= 8'hFF;
            14'h2B38: rddata <= 8'hFF; 14'h2B39: rddata <= 8'hFF; 14'h2B3A: rddata <= 8'hFF; 14'h2B3B: rddata <= 8'hFF;
            14'h2B3C: rddata <= 8'hFF; 14'h2B3D: rddata <= 8'hFF; 14'h2B3E: rddata <= 8'hFF; 14'h2B3F: rddata <= 8'hFF;
            14'h2B40: rddata <= 8'hFF; 14'h2B41: rddata <= 8'hFF; 14'h2B42: rddata <= 8'hFF; 14'h2B43: rddata <= 8'hFF;
            14'h2B44: rddata <= 8'hFF; 14'h2B45: rddata <= 8'hFF; 14'h2B46: rddata <= 8'hFF; 14'h2B47: rddata <= 8'hFF;
            14'h2B48: rddata <= 8'hFF; 14'h2B49: rddata <= 8'hFF; 14'h2B4A: rddata <= 8'hFF; 14'h2B4B: rddata <= 8'hFF;
            14'h2B4C: rddata <= 8'hFF; 14'h2B4D: rddata <= 8'hFF; 14'h2B4E: rddata <= 8'hFF; 14'h2B4F: rddata <= 8'hFF;
            14'h2B50: rddata <= 8'hFF; 14'h2B51: rddata <= 8'hFF; 14'h2B52: rddata <= 8'hFF; 14'h2B53: rddata <= 8'hFF;
            14'h2B54: rddata <= 8'hFF; 14'h2B55: rddata <= 8'hFF; 14'h2B56: rddata <= 8'hFF; 14'h2B57: rddata <= 8'hFF;
            14'h2B58: rddata <= 8'hFF; 14'h2B59: rddata <= 8'hFF; 14'h2B5A: rddata <= 8'hFF; 14'h2B5B: rddata <= 8'hFF;
            14'h2B5C: rddata <= 8'hFF; 14'h2B5D: rddata <= 8'hFF; 14'h2B5E: rddata <= 8'hFF; 14'h2B5F: rddata <= 8'hFF;
            14'h2B60: rddata <= 8'hFF; 14'h2B61: rddata <= 8'hFF; 14'h2B62: rddata <= 8'hFF; 14'h2B63: rddata <= 8'hFF;
            14'h2B64: rddata <= 8'hFF; 14'h2B65: rddata <= 8'hFF; 14'h2B66: rddata <= 8'hFF; 14'h2B67: rddata <= 8'hFF;
            14'h2B68: rddata <= 8'hFF; 14'h2B69: rddata <= 8'hFF; 14'h2B6A: rddata <= 8'hFF; 14'h2B6B: rddata <= 8'hFF;
            14'h2B6C: rddata <= 8'hFF; 14'h2B6D: rddata <= 8'hFF; 14'h2B6E: rddata <= 8'hFF; 14'h2B6F: rddata <= 8'hFF;
            14'h2B70: rddata <= 8'hFF; 14'h2B71: rddata <= 8'hFF; 14'h2B72: rddata <= 8'hFF; 14'h2B73: rddata <= 8'hFF;
            14'h2B74: rddata <= 8'hFF; 14'h2B75: rddata <= 8'hFF; 14'h2B76: rddata <= 8'hFF; 14'h2B77: rddata <= 8'hFF;
            14'h2B78: rddata <= 8'hFF; 14'h2B79: rddata <= 8'hFF; 14'h2B7A: rddata <= 8'hFF; 14'h2B7B: rddata <= 8'hFF;
            14'h2B7C: rddata <= 8'hFF; 14'h2B7D: rddata <= 8'hFF; 14'h2B7E: rddata <= 8'hFF; 14'h2B7F: rddata <= 8'hFF;
            14'h2B80: rddata <= 8'hFF; 14'h2B81: rddata <= 8'hFF; 14'h2B82: rddata <= 8'hFF; 14'h2B83: rddata <= 8'hFF;
            14'h2B84: rddata <= 8'hFF; 14'h2B85: rddata <= 8'hFF; 14'h2B86: rddata <= 8'hFF; 14'h2B87: rddata <= 8'hFF;
            14'h2B88: rddata <= 8'hFF; 14'h2B89: rddata <= 8'hFF; 14'h2B8A: rddata <= 8'hFF; 14'h2B8B: rddata <= 8'hFF;
            14'h2B8C: rddata <= 8'hFF; 14'h2B8D: rddata <= 8'hFF; 14'h2B8E: rddata <= 8'hFF; 14'h2B8F: rddata <= 8'hFF;
            14'h2B90: rddata <= 8'hFF; 14'h2B91: rddata <= 8'hFF; 14'h2B92: rddata <= 8'hFF; 14'h2B93: rddata <= 8'hFF;
            14'h2B94: rddata <= 8'hFF; 14'h2B95: rddata <= 8'hFF; 14'h2B96: rddata <= 8'hFF; 14'h2B97: rddata <= 8'hFF;
            14'h2B98: rddata <= 8'hFF; 14'h2B99: rddata <= 8'hFF; 14'h2B9A: rddata <= 8'hFF; 14'h2B9B: rddata <= 8'hFF;
            14'h2B9C: rddata <= 8'hFF; 14'h2B9D: rddata <= 8'hFF; 14'h2B9E: rddata <= 8'hFF; 14'h2B9F: rddata <= 8'hFF;
            14'h2BA0: rddata <= 8'hFF; 14'h2BA1: rddata <= 8'hFF; 14'h2BA2: rddata <= 8'hFF; 14'h2BA3: rddata <= 8'hFF;
            14'h2BA4: rddata <= 8'hFF; 14'h2BA5: rddata <= 8'hFF; 14'h2BA6: rddata <= 8'hFF; 14'h2BA7: rddata <= 8'hFF;
            14'h2BA8: rddata <= 8'hFF; 14'h2BA9: rddata <= 8'hFF; 14'h2BAA: rddata <= 8'hFF; 14'h2BAB: rddata <= 8'hFF;
            14'h2BAC: rddata <= 8'hFF; 14'h2BAD: rddata <= 8'hFF; 14'h2BAE: rddata <= 8'hFF; 14'h2BAF: rddata <= 8'hFF;
            14'h2BB0: rddata <= 8'hFF; 14'h2BB1: rddata <= 8'hFF; 14'h2BB2: rddata <= 8'hFF; 14'h2BB3: rddata <= 8'hFF;
            14'h2BB4: rddata <= 8'hFF; 14'h2BB5: rddata <= 8'hFF; 14'h2BB6: rddata <= 8'hFF; 14'h2BB7: rddata <= 8'hFF;
            14'h2BB8: rddata <= 8'hFF; 14'h2BB9: rddata <= 8'hFF; 14'h2BBA: rddata <= 8'hFF; 14'h2BBB: rddata <= 8'hFF;
            14'h2BBC: rddata <= 8'hFF; 14'h2BBD: rddata <= 8'hFF; 14'h2BBE: rddata <= 8'hFF; 14'h2BBF: rddata <= 8'hFF;
            14'h2BC0: rddata <= 8'hFF; 14'h2BC1: rddata <= 8'hFF; 14'h2BC2: rddata <= 8'hFF; 14'h2BC3: rddata <= 8'hFF;
            14'h2BC4: rddata <= 8'hFF; 14'h2BC5: rddata <= 8'hFF; 14'h2BC6: rddata <= 8'hFF; 14'h2BC7: rddata <= 8'hFF;
            14'h2BC8: rddata <= 8'hFF; 14'h2BC9: rddata <= 8'hFF; 14'h2BCA: rddata <= 8'hFF; 14'h2BCB: rddata <= 8'hFF;
            14'h2BCC: rddata <= 8'hFF; 14'h2BCD: rddata <= 8'hFF; 14'h2BCE: rddata <= 8'hFF; 14'h2BCF: rddata <= 8'hFF;
            14'h2BD0: rddata <= 8'hFF; 14'h2BD1: rddata <= 8'hFF; 14'h2BD2: rddata <= 8'hFF; 14'h2BD3: rddata <= 8'hFF;
            14'h2BD4: rddata <= 8'hFF; 14'h2BD5: rddata <= 8'hFF; 14'h2BD6: rddata <= 8'hFF; 14'h2BD7: rddata <= 8'hFF;
            14'h2BD8: rddata <= 8'hFF; 14'h2BD9: rddata <= 8'hFF; 14'h2BDA: rddata <= 8'hFF; 14'h2BDB: rddata <= 8'hFF;
            14'h2BDC: rddata <= 8'hFF; 14'h2BDD: rddata <= 8'hFF; 14'h2BDE: rddata <= 8'hFF; 14'h2BDF: rddata <= 8'hFF;
            14'h2BE0: rddata <= 8'hFF; 14'h2BE1: rddata <= 8'hFF; 14'h2BE2: rddata <= 8'hFF; 14'h2BE3: rddata <= 8'hFF;
            14'h2BE4: rddata <= 8'hFF; 14'h2BE5: rddata <= 8'hFF; 14'h2BE6: rddata <= 8'hFF; 14'h2BE7: rddata <= 8'hFF;
            14'h2BE8: rddata <= 8'hFF; 14'h2BE9: rddata <= 8'hFF; 14'h2BEA: rddata <= 8'hFF; 14'h2BEB: rddata <= 8'hFF;
            14'h2BEC: rddata <= 8'hFF; 14'h2BED: rddata <= 8'hFF; 14'h2BEE: rddata <= 8'hFF; 14'h2BEF: rddata <= 8'hFF;
            14'h2BF0: rddata <= 8'hFF; 14'h2BF1: rddata <= 8'hFF; 14'h2BF2: rddata <= 8'hFF; 14'h2BF3: rddata <= 8'hFF;
            14'h2BF4: rddata <= 8'hFF; 14'h2BF5: rddata <= 8'hFF; 14'h2BF6: rddata <= 8'hFF; 14'h2BF7: rddata <= 8'hFF;
            14'h2BF8: rddata <= 8'hFF; 14'h2BF9: rddata <= 8'hFF; 14'h2BFA: rddata <= 8'hFF; 14'h2BFB: rddata <= 8'hFF;
            14'h2BFC: rddata <= 8'hFF; 14'h2BFD: rddata <= 8'hFF; 14'h2BFE: rddata <= 8'hFF; 14'h2BFF: rddata <= 8'hFF;
            14'h2C00: rddata <= 8'hFF; 14'h2C01: rddata <= 8'hFF; 14'h2C02: rddata <= 8'hFF; 14'h2C03: rddata <= 8'hFF;
            14'h2C04: rddata <= 8'hFF; 14'h2C05: rddata <= 8'hFF; 14'h2C06: rddata <= 8'hFF; 14'h2C07: rddata <= 8'hFF;
            14'h2C08: rddata <= 8'hFF; 14'h2C09: rddata <= 8'hFF; 14'h2C0A: rddata <= 8'hFF; 14'h2C0B: rddata <= 8'hFF;
            14'h2C0C: rddata <= 8'hFF; 14'h2C0D: rddata <= 8'hFF; 14'h2C0E: rddata <= 8'hFF; 14'h2C0F: rddata <= 8'hFF;
            14'h2C10: rddata <= 8'hFF; 14'h2C11: rddata <= 8'hFF; 14'h2C12: rddata <= 8'hFF; 14'h2C13: rddata <= 8'hFF;
            14'h2C14: rddata <= 8'hFF; 14'h2C15: rddata <= 8'hFF; 14'h2C16: rddata <= 8'hFF; 14'h2C17: rddata <= 8'hFF;
            14'h2C18: rddata <= 8'hFF; 14'h2C19: rddata <= 8'hFF; 14'h2C1A: rddata <= 8'hFF; 14'h2C1B: rddata <= 8'hFF;
            14'h2C1C: rddata <= 8'hFF; 14'h2C1D: rddata <= 8'hFF; 14'h2C1E: rddata <= 8'hFF; 14'h2C1F: rddata <= 8'hFF;
            14'h2C20: rddata <= 8'hFF; 14'h2C21: rddata <= 8'hFF; 14'h2C22: rddata <= 8'hFF; 14'h2C23: rddata <= 8'hFF;
            14'h2C24: rddata <= 8'hFF; 14'h2C25: rddata <= 8'hFF; 14'h2C26: rddata <= 8'hFF; 14'h2C27: rddata <= 8'hFF;
            14'h2C28: rddata <= 8'hFF; 14'h2C29: rddata <= 8'hFF; 14'h2C2A: rddata <= 8'hFF; 14'h2C2B: rddata <= 8'hFF;
            14'h2C2C: rddata <= 8'hFF; 14'h2C2D: rddata <= 8'hFF; 14'h2C2E: rddata <= 8'hFF; 14'h2C2F: rddata <= 8'hFF;
            14'h2C30: rddata <= 8'hFF; 14'h2C31: rddata <= 8'hFF; 14'h2C32: rddata <= 8'hFF; 14'h2C33: rddata <= 8'hFF;
            14'h2C34: rddata <= 8'hFF; 14'h2C35: rddata <= 8'hFF; 14'h2C36: rddata <= 8'hFF; 14'h2C37: rddata <= 8'hFF;
            14'h2C38: rddata <= 8'hFF; 14'h2C39: rddata <= 8'hFF; 14'h2C3A: rddata <= 8'hFF; 14'h2C3B: rddata <= 8'hFF;
            14'h2C3C: rddata <= 8'hFF; 14'h2C3D: rddata <= 8'hFF; 14'h2C3E: rddata <= 8'hFF; 14'h2C3F: rddata <= 8'hFF;
            14'h2C40: rddata <= 8'hFF; 14'h2C41: rddata <= 8'hFF; 14'h2C42: rddata <= 8'hFF; 14'h2C43: rddata <= 8'hFF;
            14'h2C44: rddata <= 8'hFF; 14'h2C45: rddata <= 8'hFF; 14'h2C46: rddata <= 8'hFF; 14'h2C47: rddata <= 8'hFF;
            14'h2C48: rddata <= 8'hFF; 14'h2C49: rddata <= 8'hFF; 14'h2C4A: rddata <= 8'hFF; 14'h2C4B: rddata <= 8'hFF;
            14'h2C4C: rddata <= 8'hFF; 14'h2C4D: rddata <= 8'hFF; 14'h2C4E: rddata <= 8'hFF; 14'h2C4F: rddata <= 8'hFF;
            14'h2C50: rddata <= 8'hFF; 14'h2C51: rddata <= 8'hFF; 14'h2C52: rddata <= 8'hFF; 14'h2C53: rddata <= 8'hFF;
            14'h2C54: rddata <= 8'hFF; 14'h2C55: rddata <= 8'hFF; 14'h2C56: rddata <= 8'hFF; 14'h2C57: rddata <= 8'hFF;
            14'h2C58: rddata <= 8'hFF; 14'h2C59: rddata <= 8'hFF; 14'h2C5A: rddata <= 8'hFF; 14'h2C5B: rddata <= 8'hFF;
            14'h2C5C: rddata <= 8'hFF; 14'h2C5D: rddata <= 8'hFF; 14'h2C5E: rddata <= 8'hFF; 14'h2C5F: rddata <= 8'hFF;
            14'h2C60: rddata <= 8'hFF; 14'h2C61: rddata <= 8'hFF; 14'h2C62: rddata <= 8'hFF; 14'h2C63: rddata <= 8'hFF;
            14'h2C64: rddata <= 8'hFF; 14'h2C65: rddata <= 8'hFF; 14'h2C66: rddata <= 8'hFF; 14'h2C67: rddata <= 8'hFF;
            14'h2C68: rddata <= 8'hFF; 14'h2C69: rddata <= 8'hFF; 14'h2C6A: rddata <= 8'hFF; 14'h2C6B: rddata <= 8'hFF;
            14'h2C6C: rddata <= 8'hFF; 14'h2C6D: rddata <= 8'hFF; 14'h2C6E: rddata <= 8'hFF; 14'h2C6F: rddata <= 8'hFF;
            14'h2C70: rddata <= 8'hFF; 14'h2C71: rddata <= 8'hFF; 14'h2C72: rddata <= 8'hFF; 14'h2C73: rddata <= 8'hFF;
            14'h2C74: rddata <= 8'hFF; 14'h2C75: rddata <= 8'hFF; 14'h2C76: rddata <= 8'hFF; 14'h2C77: rddata <= 8'hFF;
            14'h2C78: rddata <= 8'hFF; 14'h2C79: rddata <= 8'hFF; 14'h2C7A: rddata <= 8'hFF; 14'h2C7B: rddata <= 8'hFF;
            14'h2C7C: rddata <= 8'hFF; 14'h2C7D: rddata <= 8'hFF; 14'h2C7E: rddata <= 8'hFF; 14'h2C7F: rddata <= 8'hFF;
            14'h2C80: rddata <= 8'hFF; 14'h2C81: rddata <= 8'hFF; 14'h2C82: rddata <= 8'hFF; 14'h2C83: rddata <= 8'hFF;
            14'h2C84: rddata <= 8'hFF; 14'h2C85: rddata <= 8'hFF; 14'h2C86: rddata <= 8'hFF; 14'h2C87: rddata <= 8'hFF;
            14'h2C88: rddata <= 8'hFF; 14'h2C89: rddata <= 8'hFF; 14'h2C8A: rddata <= 8'hFF; 14'h2C8B: rddata <= 8'hFF;
            14'h2C8C: rddata <= 8'hFF; 14'h2C8D: rddata <= 8'hFF; 14'h2C8E: rddata <= 8'hFF; 14'h2C8F: rddata <= 8'hFF;
            14'h2C90: rddata <= 8'hFF; 14'h2C91: rddata <= 8'hFF; 14'h2C92: rddata <= 8'hFF; 14'h2C93: rddata <= 8'hFF;
            14'h2C94: rddata <= 8'hFF; 14'h2C95: rddata <= 8'hFF; 14'h2C96: rddata <= 8'hFF; 14'h2C97: rddata <= 8'hFF;
            14'h2C98: rddata <= 8'hFF; 14'h2C99: rddata <= 8'hFF; 14'h2C9A: rddata <= 8'hFF; 14'h2C9B: rddata <= 8'hFF;
            14'h2C9C: rddata <= 8'hFF; 14'h2C9D: rddata <= 8'hFF; 14'h2C9E: rddata <= 8'hFF; 14'h2C9F: rddata <= 8'hFF;
            14'h2CA0: rddata <= 8'hFF; 14'h2CA1: rddata <= 8'hFF; 14'h2CA2: rddata <= 8'hFF; 14'h2CA3: rddata <= 8'hFF;
            14'h2CA4: rddata <= 8'hFF; 14'h2CA5: rddata <= 8'hFF; 14'h2CA6: rddata <= 8'hFF; 14'h2CA7: rddata <= 8'hFF;
            14'h2CA8: rddata <= 8'hFF; 14'h2CA9: rddata <= 8'hFF; 14'h2CAA: rddata <= 8'hFF; 14'h2CAB: rddata <= 8'hFF;
            14'h2CAC: rddata <= 8'hFF; 14'h2CAD: rddata <= 8'hFF; 14'h2CAE: rddata <= 8'hFF; 14'h2CAF: rddata <= 8'hFF;
            14'h2CB0: rddata <= 8'hFF; 14'h2CB1: rddata <= 8'hFF; 14'h2CB2: rddata <= 8'hFF; 14'h2CB3: rddata <= 8'hFF;
            14'h2CB4: rddata <= 8'hFF; 14'h2CB5: rddata <= 8'hFF; 14'h2CB6: rddata <= 8'hFF; 14'h2CB7: rddata <= 8'hFF;
            14'h2CB8: rddata <= 8'hFF; 14'h2CB9: rddata <= 8'hFF; 14'h2CBA: rddata <= 8'hFF; 14'h2CBB: rddata <= 8'hFF;
            14'h2CBC: rddata <= 8'hFF; 14'h2CBD: rddata <= 8'hFF; 14'h2CBE: rddata <= 8'hFF; 14'h2CBF: rddata <= 8'hFF;
            14'h2CC0: rddata <= 8'hFF; 14'h2CC1: rddata <= 8'hFF; 14'h2CC2: rddata <= 8'hFF; 14'h2CC3: rddata <= 8'hFF;
            14'h2CC4: rddata <= 8'hFF; 14'h2CC5: rddata <= 8'hFF; 14'h2CC6: rddata <= 8'hFF; 14'h2CC7: rddata <= 8'hFF;
            14'h2CC8: rddata <= 8'hFF; 14'h2CC9: rddata <= 8'hFF; 14'h2CCA: rddata <= 8'hFF; 14'h2CCB: rddata <= 8'hFF;
            14'h2CCC: rddata <= 8'hFF; 14'h2CCD: rddata <= 8'hFF; 14'h2CCE: rddata <= 8'hFF; 14'h2CCF: rddata <= 8'hFF;
            14'h2CD0: rddata <= 8'hFF; 14'h2CD1: rddata <= 8'hFF; 14'h2CD2: rddata <= 8'hFF; 14'h2CD3: rddata <= 8'hFF;
            14'h2CD4: rddata <= 8'hFF; 14'h2CD5: rddata <= 8'hFF; 14'h2CD6: rddata <= 8'hFF; 14'h2CD7: rddata <= 8'hFF;
            14'h2CD8: rddata <= 8'hFF; 14'h2CD9: rddata <= 8'hFF; 14'h2CDA: rddata <= 8'hFF; 14'h2CDB: rddata <= 8'hFF;
            14'h2CDC: rddata <= 8'hFF; 14'h2CDD: rddata <= 8'hFF; 14'h2CDE: rddata <= 8'hFF; 14'h2CDF: rddata <= 8'hFF;
            14'h2CE0: rddata <= 8'hFF; 14'h2CE1: rddata <= 8'hFF; 14'h2CE2: rddata <= 8'hFF; 14'h2CE3: rddata <= 8'hFF;
            14'h2CE4: rddata <= 8'hFF; 14'h2CE5: rddata <= 8'hFF; 14'h2CE6: rddata <= 8'hFF; 14'h2CE7: rddata <= 8'hFF;
            14'h2CE8: rddata <= 8'hFF; 14'h2CE9: rddata <= 8'hFF; 14'h2CEA: rddata <= 8'hFF; 14'h2CEB: rddata <= 8'hFF;
            14'h2CEC: rddata <= 8'hFF; 14'h2CED: rddata <= 8'hFF; 14'h2CEE: rddata <= 8'hFF; 14'h2CEF: rddata <= 8'hFF;
            14'h2CF0: rddata <= 8'hFF; 14'h2CF1: rddata <= 8'hFF; 14'h2CF2: rddata <= 8'hFF; 14'h2CF3: rddata <= 8'hFF;
            14'h2CF4: rddata <= 8'hFF; 14'h2CF5: rddata <= 8'hFF; 14'h2CF6: rddata <= 8'hFF; 14'h2CF7: rddata <= 8'hFF;
            14'h2CF8: rddata <= 8'hFF; 14'h2CF9: rddata <= 8'hFF; 14'h2CFA: rddata <= 8'hFF; 14'h2CFB: rddata <= 8'hFF;
            14'h2CFC: rddata <= 8'hFF; 14'h2CFD: rddata <= 8'hFF; 14'h2CFE: rddata <= 8'hFF; 14'h2CFF: rddata <= 8'hFF;
            14'h2D00: rddata <= 8'hFF; 14'h2D01: rddata <= 8'hFF; 14'h2D02: rddata <= 8'hFF; 14'h2D03: rddata <= 8'hFF;
            14'h2D04: rddata <= 8'hFF; 14'h2D05: rddata <= 8'hFF; 14'h2D06: rddata <= 8'hFF; 14'h2D07: rddata <= 8'hFF;
            14'h2D08: rddata <= 8'hFF; 14'h2D09: rddata <= 8'hFF; 14'h2D0A: rddata <= 8'hFF; 14'h2D0B: rddata <= 8'hFF;
            14'h2D0C: rddata <= 8'hFF; 14'h2D0D: rddata <= 8'hFF; 14'h2D0E: rddata <= 8'hFF; 14'h2D0F: rddata <= 8'hFF;
            14'h2D10: rddata <= 8'hFF; 14'h2D11: rddata <= 8'hFF; 14'h2D12: rddata <= 8'hFF; 14'h2D13: rddata <= 8'hFF;
            14'h2D14: rddata <= 8'hFF; 14'h2D15: rddata <= 8'hFF; 14'h2D16: rddata <= 8'hFF; 14'h2D17: rddata <= 8'hFF;
            14'h2D18: rddata <= 8'hFF; 14'h2D19: rddata <= 8'hFF; 14'h2D1A: rddata <= 8'hFF; 14'h2D1B: rddata <= 8'hFF;
            14'h2D1C: rddata <= 8'hFF; 14'h2D1D: rddata <= 8'hFF; 14'h2D1E: rddata <= 8'hFF; 14'h2D1F: rddata <= 8'hFF;
            14'h2D20: rddata <= 8'hFF; 14'h2D21: rddata <= 8'hFF; 14'h2D22: rddata <= 8'hFF; 14'h2D23: rddata <= 8'hFF;
            14'h2D24: rddata <= 8'hFF; 14'h2D25: rddata <= 8'hFF; 14'h2D26: rddata <= 8'hFF; 14'h2D27: rddata <= 8'hFF;
            14'h2D28: rddata <= 8'hFF; 14'h2D29: rddata <= 8'hFF; 14'h2D2A: rddata <= 8'hFF; 14'h2D2B: rddata <= 8'hFF;
            14'h2D2C: rddata <= 8'hFF; 14'h2D2D: rddata <= 8'hFF; 14'h2D2E: rddata <= 8'hFF; 14'h2D2F: rddata <= 8'hFF;
            14'h2D30: rddata <= 8'hFF; 14'h2D31: rddata <= 8'hFF; 14'h2D32: rddata <= 8'hFF; 14'h2D33: rddata <= 8'hFF;
            14'h2D34: rddata <= 8'hFF; 14'h2D35: rddata <= 8'hFF; 14'h2D36: rddata <= 8'hFF; 14'h2D37: rddata <= 8'hFF;
            14'h2D38: rddata <= 8'hFF; 14'h2D39: rddata <= 8'hFF; 14'h2D3A: rddata <= 8'hFF; 14'h2D3B: rddata <= 8'hFF;
            14'h2D3C: rddata <= 8'hFF; 14'h2D3D: rddata <= 8'hFF; 14'h2D3E: rddata <= 8'hFF; 14'h2D3F: rddata <= 8'hFF;
            14'h2D40: rddata <= 8'hFF; 14'h2D41: rddata <= 8'hFF; 14'h2D42: rddata <= 8'hFF; 14'h2D43: rddata <= 8'hFF;
            14'h2D44: rddata <= 8'hFF; 14'h2D45: rddata <= 8'hFF; 14'h2D46: rddata <= 8'hFF; 14'h2D47: rddata <= 8'hFF;
            14'h2D48: rddata <= 8'hFF; 14'h2D49: rddata <= 8'hFF; 14'h2D4A: rddata <= 8'hFF; 14'h2D4B: rddata <= 8'hFF;
            14'h2D4C: rddata <= 8'hFF; 14'h2D4D: rddata <= 8'hFF; 14'h2D4E: rddata <= 8'hFF; 14'h2D4F: rddata <= 8'hFF;
            14'h2D50: rddata <= 8'hFF; 14'h2D51: rddata <= 8'hFF; 14'h2D52: rddata <= 8'hFF; 14'h2D53: rddata <= 8'hFF;
            14'h2D54: rddata <= 8'hFF; 14'h2D55: rddata <= 8'hFF; 14'h2D56: rddata <= 8'hFF; 14'h2D57: rddata <= 8'hFF;
            14'h2D58: rddata <= 8'hFF; 14'h2D59: rddata <= 8'hFF; 14'h2D5A: rddata <= 8'hFF; 14'h2D5B: rddata <= 8'hFF;
            14'h2D5C: rddata <= 8'hFF; 14'h2D5D: rddata <= 8'hFF; 14'h2D5E: rddata <= 8'hFF; 14'h2D5F: rddata <= 8'hFF;
            14'h2D60: rddata <= 8'hFF; 14'h2D61: rddata <= 8'hFF; 14'h2D62: rddata <= 8'hFF; 14'h2D63: rddata <= 8'hFF;
            14'h2D64: rddata <= 8'hFF; 14'h2D65: rddata <= 8'hFF; 14'h2D66: rddata <= 8'hFF; 14'h2D67: rddata <= 8'hFF;
            14'h2D68: rddata <= 8'hFF; 14'h2D69: rddata <= 8'hFF; 14'h2D6A: rddata <= 8'hFF; 14'h2D6B: rddata <= 8'hFF;
            14'h2D6C: rddata <= 8'hFF; 14'h2D6D: rddata <= 8'hFF; 14'h2D6E: rddata <= 8'hFF; 14'h2D6F: rddata <= 8'hFF;
            14'h2D70: rddata <= 8'hFF; 14'h2D71: rddata <= 8'hFF; 14'h2D72: rddata <= 8'hFF; 14'h2D73: rddata <= 8'hFF;
            14'h2D74: rddata <= 8'hFF; 14'h2D75: rddata <= 8'hFF; 14'h2D76: rddata <= 8'hFF; 14'h2D77: rddata <= 8'hFF;
            14'h2D78: rddata <= 8'hFF; 14'h2D79: rddata <= 8'hFF; 14'h2D7A: rddata <= 8'hFF; 14'h2D7B: rddata <= 8'hFF;
            14'h2D7C: rddata <= 8'hFF; 14'h2D7D: rddata <= 8'hFF; 14'h2D7E: rddata <= 8'hFF; 14'h2D7F: rddata <= 8'hFF;
            14'h2D80: rddata <= 8'hFF; 14'h2D81: rddata <= 8'hFF; 14'h2D82: rddata <= 8'hFF; 14'h2D83: rddata <= 8'hFF;
            14'h2D84: rddata <= 8'hFF; 14'h2D85: rddata <= 8'hFF; 14'h2D86: rddata <= 8'hFF; 14'h2D87: rddata <= 8'hFF;
            14'h2D88: rddata <= 8'hFF; 14'h2D89: rddata <= 8'hFF; 14'h2D8A: rddata <= 8'hFF; 14'h2D8B: rddata <= 8'hFF;
            14'h2D8C: rddata <= 8'hFF; 14'h2D8D: rddata <= 8'hFF; 14'h2D8E: rddata <= 8'hFF; 14'h2D8F: rddata <= 8'hFF;
            14'h2D90: rddata <= 8'hFF; 14'h2D91: rddata <= 8'hFF; 14'h2D92: rddata <= 8'hFF; 14'h2D93: rddata <= 8'hFF;
            14'h2D94: rddata <= 8'hFF; 14'h2D95: rddata <= 8'hFF; 14'h2D96: rddata <= 8'hFF; 14'h2D97: rddata <= 8'hFF;
            14'h2D98: rddata <= 8'hFF; 14'h2D99: rddata <= 8'hFF; 14'h2D9A: rddata <= 8'hFF; 14'h2D9B: rddata <= 8'hFF;
            14'h2D9C: rddata <= 8'hFF; 14'h2D9D: rddata <= 8'hFF; 14'h2D9E: rddata <= 8'hFF; 14'h2D9F: rddata <= 8'hFF;
            14'h2DA0: rddata <= 8'hFF; 14'h2DA1: rddata <= 8'hFF; 14'h2DA2: rddata <= 8'hFF; 14'h2DA3: rddata <= 8'hFF;
            14'h2DA4: rddata <= 8'hFF; 14'h2DA5: rddata <= 8'hFF; 14'h2DA6: rddata <= 8'hFF; 14'h2DA7: rddata <= 8'hFF;
            14'h2DA8: rddata <= 8'hFF; 14'h2DA9: rddata <= 8'hFF; 14'h2DAA: rddata <= 8'hFF; 14'h2DAB: rddata <= 8'hFF;
            14'h2DAC: rddata <= 8'hFF; 14'h2DAD: rddata <= 8'hFF; 14'h2DAE: rddata <= 8'hFF; 14'h2DAF: rddata <= 8'hFF;
            14'h2DB0: rddata <= 8'hFF; 14'h2DB1: rddata <= 8'hFF; 14'h2DB2: rddata <= 8'hFF; 14'h2DB3: rddata <= 8'hFF;
            14'h2DB4: rddata <= 8'hFF; 14'h2DB5: rddata <= 8'hFF; 14'h2DB6: rddata <= 8'hFF; 14'h2DB7: rddata <= 8'hFF;
            14'h2DB8: rddata <= 8'hFF; 14'h2DB9: rddata <= 8'hFF; 14'h2DBA: rddata <= 8'hFF; 14'h2DBB: rddata <= 8'hFF;
            14'h2DBC: rddata <= 8'hFF; 14'h2DBD: rddata <= 8'hFF; 14'h2DBE: rddata <= 8'hFF; 14'h2DBF: rddata <= 8'hFF;
            14'h2DC0: rddata <= 8'hFF; 14'h2DC1: rddata <= 8'hFF; 14'h2DC2: rddata <= 8'hFF; 14'h2DC3: rddata <= 8'hFF;
            14'h2DC4: rddata <= 8'hFF; 14'h2DC5: rddata <= 8'hFF; 14'h2DC6: rddata <= 8'hFF; 14'h2DC7: rddata <= 8'hFF;
            14'h2DC8: rddata <= 8'hFF; 14'h2DC9: rddata <= 8'hFF; 14'h2DCA: rddata <= 8'hFF; 14'h2DCB: rddata <= 8'hFF;
            14'h2DCC: rddata <= 8'hFF; 14'h2DCD: rddata <= 8'hFF; 14'h2DCE: rddata <= 8'hFF; 14'h2DCF: rddata <= 8'hFF;
            14'h2DD0: rddata <= 8'hFF; 14'h2DD1: rddata <= 8'hFF; 14'h2DD2: rddata <= 8'hFF; 14'h2DD3: rddata <= 8'hFF;
            14'h2DD4: rddata <= 8'hFF; 14'h2DD5: rddata <= 8'hFF; 14'h2DD6: rddata <= 8'hFF; 14'h2DD7: rddata <= 8'hFF;
            14'h2DD8: rddata <= 8'hFF; 14'h2DD9: rddata <= 8'hFF; 14'h2DDA: rddata <= 8'hFF; 14'h2DDB: rddata <= 8'hFF;
            14'h2DDC: rddata <= 8'hFF; 14'h2DDD: rddata <= 8'hFF; 14'h2DDE: rddata <= 8'hFF; 14'h2DDF: rddata <= 8'hFF;
            14'h2DE0: rddata <= 8'hFF; 14'h2DE1: rddata <= 8'hFF; 14'h2DE2: rddata <= 8'hFF; 14'h2DE3: rddata <= 8'hFF;
            14'h2DE4: rddata <= 8'hFF; 14'h2DE5: rddata <= 8'hFF; 14'h2DE6: rddata <= 8'hFF; 14'h2DE7: rddata <= 8'hFF;
            14'h2DE8: rddata <= 8'hFF; 14'h2DE9: rddata <= 8'hFF; 14'h2DEA: rddata <= 8'hFF; 14'h2DEB: rddata <= 8'hFF;
            14'h2DEC: rddata <= 8'hFF; 14'h2DED: rddata <= 8'hFF; 14'h2DEE: rddata <= 8'hFF; 14'h2DEF: rddata <= 8'hFF;
            14'h2DF0: rddata <= 8'hFF; 14'h2DF1: rddata <= 8'hFF; 14'h2DF2: rddata <= 8'hFF; 14'h2DF3: rddata <= 8'hFF;
            14'h2DF4: rddata <= 8'hFF; 14'h2DF5: rddata <= 8'hFF; 14'h2DF6: rddata <= 8'hFF; 14'h2DF7: rddata <= 8'hFF;
            14'h2DF8: rddata <= 8'hFF; 14'h2DF9: rddata <= 8'hFF; 14'h2DFA: rddata <= 8'hFF; 14'h2DFB: rddata <= 8'hFF;
            14'h2DFC: rddata <= 8'hFF; 14'h2DFD: rddata <= 8'hFF; 14'h2DFE: rddata <= 8'hFF; 14'h2DFF: rddata <= 8'hFF;
            14'h2E00: rddata <= 8'hFF; 14'h2E01: rddata <= 8'hFF; 14'h2E02: rddata <= 8'hFF; 14'h2E03: rddata <= 8'hFF;
            14'h2E04: rddata <= 8'hFF; 14'h2E05: rddata <= 8'hFF; 14'h2E06: rddata <= 8'hFF; 14'h2E07: rddata <= 8'hFF;
            14'h2E08: rddata <= 8'hFF; 14'h2E09: rddata <= 8'hFF; 14'h2E0A: rddata <= 8'hFF; 14'h2E0B: rddata <= 8'hFF;
            14'h2E0C: rddata <= 8'hFF; 14'h2E0D: rddata <= 8'hFF; 14'h2E0E: rddata <= 8'hFF; 14'h2E0F: rddata <= 8'hFF;
            14'h2E10: rddata <= 8'hFF; 14'h2E11: rddata <= 8'hFF; 14'h2E12: rddata <= 8'hFF; 14'h2E13: rddata <= 8'hFF;
            14'h2E14: rddata <= 8'hFF; 14'h2E15: rddata <= 8'hFF; 14'h2E16: rddata <= 8'hFF; 14'h2E17: rddata <= 8'hFF;
            14'h2E18: rddata <= 8'hFF; 14'h2E19: rddata <= 8'hFF; 14'h2E1A: rddata <= 8'hFF; 14'h2E1B: rddata <= 8'hFF;
            14'h2E1C: rddata <= 8'hFF; 14'h2E1D: rddata <= 8'hFF; 14'h2E1E: rddata <= 8'hFF; 14'h2E1F: rddata <= 8'hFF;
            14'h2E20: rddata <= 8'hFF; 14'h2E21: rddata <= 8'hFF; 14'h2E22: rddata <= 8'hFF; 14'h2E23: rddata <= 8'hFF;
            14'h2E24: rddata <= 8'hFF; 14'h2E25: rddata <= 8'hFF; 14'h2E26: rddata <= 8'hFF; 14'h2E27: rddata <= 8'hFF;
            14'h2E28: rddata <= 8'hFF; 14'h2E29: rddata <= 8'hFF; 14'h2E2A: rddata <= 8'hFF; 14'h2E2B: rddata <= 8'hFF;
            14'h2E2C: rddata <= 8'hFF; 14'h2E2D: rddata <= 8'hFF; 14'h2E2E: rddata <= 8'hFF; 14'h2E2F: rddata <= 8'hFF;
            14'h2E30: rddata <= 8'hFF; 14'h2E31: rddata <= 8'hFF; 14'h2E32: rddata <= 8'hFF; 14'h2E33: rddata <= 8'hFF;
            14'h2E34: rddata <= 8'hFF; 14'h2E35: rddata <= 8'hFF; 14'h2E36: rddata <= 8'hFF; 14'h2E37: rddata <= 8'hFF;
            14'h2E38: rddata <= 8'hFF; 14'h2E39: rddata <= 8'hFF; 14'h2E3A: rddata <= 8'hFF; 14'h2E3B: rddata <= 8'hFF;
            14'h2E3C: rddata <= 8'hFF; 14'h2E3D: rddata <= 8'hFF; 14'h2E3E: rddata <= 8'hFF; 14'h2E3F: rddata <= 8'hFF;
            14'h2E40: rddata <= 8'hFF; 14'h2E41: rddata <= 8'hFF; 14'h2E42: rddata <= 8'hFF; 14'h2E43: rddata <= 8'hFF;
            14'h2E44: rddata <= 8'hFF; 14'h2E45: rddata <= 8'hFF; 14'h2E46: rddata <= 8'hFF; 14'h2E47: rddata <= 8'hFF;
            14'h2E48: rddata <= 8'hFF; 14'h2E49: rddata <= 8'hFF; 14'h2E4A: rddata <= 8'hFF; 14'h2E4B: rddata <= 8'hFF;
            14'h2E4C: rddata <= 8'hFF; 14'h2E4D: rddata <= 8'hFF; 14'h2E4E: rddata <= 8'hFF; 14'h2E4F: rddata <= 8'hFF;
            14'h2E50: rddata <= 8'hFF; 14'h2E51: rddata <= 8'hFF; 14'h2E52: rddata <= 8'hFF; 14'h2E53: rddata <= 8'hFF;
            14'h2E54: rddata <= 8'hFF; 14'h2E55: rddata <= 8'hFF; 14'h2E56: rddata <= 8'hFF; 14'h2E57: rddata <= 8'hFF;
            14'h2E58: rddata <= 8'hFF; 14'h2E59: rddata <= 8'hFF; 14'h2E5A: rddata <= 8'hFF; 14'h2E5B: rddata <= 8'hFF;
            14'h2E5C: rddata <= 8'hFF; 14'h2E5D: rddata <= 8'hFF; 14'h2E5E: rddata <= 8'hFF; 14'h2E5F: rddata <= 8'hFF;
            14'h2E60: rddata <= 8'hFF; 14'h2E61: rddata <= 8'hFF; 14'h2E62: rddata <= 8'hFF; 14'h2E63: rddata <= 8'hFF;
            14'h2E64: rddata <= 8'hFF; 14'h2E65: rddata <= 8'hFF; 14'h2E66: rddata <= 8'hFF; 14'h2E67: rddata <= 8'hFF;
            14'h2E68: rddata <= 8'hFF; 14'h2E69: rddata <= 8'hFF; 14'h2E6A: rddata <= 8'hFF; 14'h2E6B: rddata <= 8'hFF;
            14'h2E6C: rddata <= 8'hFF; 14'h2E6D: rddata <= 8'hFF; 14'h2E6E: rddata <= 8'hFF; 14'h2E6F: rddata <= 8'hFF;
            14'h2E70: rddata <= 8'hFF; 14'h2E71: rddata <= 8'hFF; 14'h2E72: rddata <= 8'hFF; 14'h2E73: rddata <= 8'hFF;
            14'h2E74: rddata <= 8'hFF; 14'h2E75: rddata <= 8'hFF; 14'h2E76: rddata <= 8'hFF; 14'h2E77: rddata <= 8'hFF;
            14'h2E78: rddata <= 8'hFF; 14'h2E79: rddata <= 8'hFF; 14'h2E7A: rddata <= 8'hFF; 14'h2E7B: rddata <= 8'hFF;
            14'h2E7C: rddata <= 8'hFF; 14'h2E7D: rddata <= 8'hFF; 14'h2E7E: rddata <= 8'hFF; 14'h2E7F: rddata <= 8'hFF;
            14'h2E80: rddata <= 8'hFF; 14'h2E81: rddata <= 8'hFF; 14'h2E82: rddata <= 8'hFF; 14'h2E83: rddata <= 8'hFF;
            14'h2E84: rddata <= 8'hFF; 14'h2E85: rddata <= 8'hFF; 14'h2E86: rddata <= 8'hFF; 14'h2E87: rddata <= 8'hFF;
            14'h2E88: rddata <= 8'hFF; 14'h2E89: rddata <= 8'hFF; 14'h2E8A: rddata <= 8'hFF; 14'h2E8B: rddata <= 8'hFF;
            14'h2E8C: rddata <= 8'hFF; 14'h2E8D: rddata <= 8'hFF; 14'h2E8E: rddata <= 8'hFF; 14'h2E8F: rddata <= 8'hFF;
            14'h2E90: rddata <= 8'hFF; 14'h2E91: rddata <= 8'hFF; 14'h2E92: rddata <= 8'hFF; 14'h2E93: rddata <= 8'hFF;
            14'h2E94: rddata <= 8'hFF; 14'h2E95: rddata <= 8'hFF; 14'h2E96: rddata <= 8'hFF; 14'h2E97: rddata <= 8'hFF;
            14'h2E98: rddata <= 8'hFF; 14'h2E99: rddata <= 8'hFF; 14'h2E9A: rddata <= 8'hFF; 14'h2E9B: rddata <= 8'hFF;
            14'h2E9C: rddata <= 8'hFF; 14'h2E9D: rddata <= 8'hFF; 14'h2E9E: rddata <= 8'hFF; 14'h2E9F: rddata <= 8'hFF;
            14'h2EA0: rddata <= 8'hFF; 14'h2EA1: rddata <= 8'hFF; 14'h2EA2: rddata <= 8'hFF; 14'h2EA3: rddata <= 8'hFF;
            14'h2EA4: rddata <= 8'hFF; 14'h2EA5: rddata <= 8'hFF; 14'h2EA6: rddata <= 8'hFF; 14'h2EA7: rddata <= 8'hFF;
            14'h2EA8: rddata <= 8'hFF; 14'h2EA9: rddata <= 8'hFF; 14'h2EAA: rddata <= 8'hFF; 14'h2EAB: rddata <= 8'hFF;
            14'h2EAC: rddata <= 8'hFF; 14'h2EAD: rddata <= 8'hFF; 14'h2EAE: rddata <= 8'hFF; 14'h2EAF: rddata <= 8'hFF;
            14'h2EB0: rddata <= 8'hFF; 14'h2EB1: rddata <= 8'hFF; 14'h2EB2: rddata <= 8'hFF; 14'h2EB3: rddata <= 8'hFF;
            14'h2EB4: rddata <= 8'hFF; 14'h2EB5: rddata <= 8'hFF; 14'h2EB6: rddata <= 8'hFF; 14'h2EB7: rddata <= 8'hFF;
            14'h2EB8: rddata <= 8'hFF; 14'h2EB9: rddata <= 8'hFF; 14'h2EBA: rddata <= 8'hFF; 14'h2EBB: rddata <= 8'hFF;
            14'h2EBC: rddata <= 8'hFF; 14'h2EBD: rddata <= 8'hFF; 14'h2EBE: rddata <= 8'hFF; 14'h2EBF: rddata <= 8'hFF;
            14'h2EC0: rddata <= 8'hFF; 14'h2EC1: rddata <= 8'hFF; 14'h2EC2: rddata <= 8'hFF; 14'h2EC3: rddata <= 8'hFF;
            14'h2EC4: rddata <= 8'hFF; 14'h2EC5: rddata <= 8'hFF; 14'h2EC6: rddata <= 8'hFF; 14'h2EC7: rddata <= 8'hFF;
            14'h2EC8: rddata <= 8'hFF; 14'h2EC9: rddata <= 8'hFF; 14'h2ECA: rddata <= 8'hFF; 14'h2ECB: rddata <= 8'hFF;
            14'h2ECC: rddata <= 8'hFF; 14'h2ECD: rddata <= 8'hFF; 14'h2ECE: rddata <= 8'hFF; 14'h2ECF: rddata <= 8'hFF;
            14'h2ED0: rddata <= 8'hFF; 14'h2ED1: rddata <= 8'hFF; 14'h2ED2: rddata <= 8'hFF; 14'h2ED3: rddata <= 8'hFF;
            14'h2ED4: rddata <= 8'hFF; 14'h2ED5: rddata <= 8'hFF; 14'h2ED6: rddata <= 8'hFF; 14'h2ED7: rddata <= 8'hFF;
            14'h2ED8: rddata <= 8'hFF; 14'h2ED9: rddata <= 8'hFF; 14'h2EDA: rddata <= 8'hFF; 14'h2EDB: rddata <= 8'hFF;
            14'h2EDC: rddata <= 8'hFF; 14'h2EDD: rddata <= 8'hFF; 14'h2EDE: rddata <= 8'hFF; 14'h2EDF: rddata <= 8'hFF;
            14'h2EE0: rddata <= 8'hFF; 14'h2EE1: rddata <= 8'hFF; 14'h2EE2: rddata <= 8'hFF; 14'h2EE3: rddata <= 8'hFF;
            14'h2EE4: rddata <= 8'hFF; 14'h2EE5: rddata <= 8'hFF; 14'h2EE6: rddata <= 8'hFF; 14'h2EE7: rddata <= 8'hFF;
            14'h2EE8: rddata <= 8'hFF; 14'h2EE9: rddata <= 8'hFF; 14'h2EEA: rddata <= 8'hFF; 14'h2EEB: rddata <= 8'hFF;
            14'h2EEC: rddata <= 8'hFF; 14'h2EED: rddata <= 8'hFF; 14'h2EEE: rddata <= 8'hFF; 14'h2EEF: rddata <= 8'hFF;
            14'h2EF0: rddata <= 8'hFF; 14'h2EF1: rddata <= 8'hFF; 14'h2EF2: rddata <= 8'hFF; 14'h2EF3: rddata <= 8'hFF;
            14'h2EF4: rddata <= 8'hFF; 14'h2EF5: rddata <= 8'hFF; 14'h2EF6: rddata <= 8'hFF; 14'h2EF7: rddata <= 8'hFF;
            14'h2EF8: rddata <= 8'hFF; 14'h2EF9: rddata <= 8'hFF; 14'h2EFA: rddata <= 8'hFF; 14'h2EFB: rddata <= 8'hFF;
            14'h2EFC: rddata <= 8'hFF; 14'h2EFD: rddata <= 8'hFF; 14'h2EFE: rddata <= 8'hFF; 14'h2EFF: rddata <= 8'hFF;
            14'h2F00: rddata <= 8'hFF; 14'h2F01: rddata <= 8'hFF; 14'h2F02: rddata <= 8'hFF; 14'h2F03: rddata <= 8'hFF;
            14'h2F04: rddata <= 8'hFF; 14'h2F05: rddata <= 8'hFF; 14'h2F06: rddata <= 8'hFF; 14'h2F07: rddata <= 8'hFF;
            14'h2F08: rddata <= 8'hFF; 14'h2F09: rddata <= 8'hFF; 14'h2F0A: rddata <= 8'hFF; 14'h2F0B: rddata <= 8'hFF;
            14'h2F0C: rddata <= 8'hFF; 14'h2F0D: rddata <= 8'hFF; 14'h2F0E: rddata <= 8'hFF; 14'h2F0F: rddata <= 8'hFF;
            14'h2F10: rddata <= 8'hFF; 14'h2F11: rddata <= 8'hFF; 14'h2F12: rddata <= 8'hFF; 14'h2F13: rddata <= 8'hFF;
            14'h2F14: rddata <= 8'hFF; 14'h2F15: rddata <= 8'hFF; 14'h2F16: rddata <= 8'hFF; 14'h2F17: rddata <= 8'hFF;
            14'h2F18: rddata <= 8'hFF; 14'h2F19: rddata <= 8'hFF; 14'h2F1A: rddata <= 8'hFF; 14'h2F1B: rddata <= 8'hFF;
            14'h2F1C: rddata <= 8'hFF; 14'h2F1D: rddata <= 8'hFF; 14'h2F1E: rddata <= 8'hFF; 14'h2F1F: rddata <= 8'hFF;
            14'h2F20: rddata <= 8'hFF; 14'h2F21: rddata <= 8'hFF; 14'h2F22: rddata <= 8'hFF; 14'h2F23: rddata <= 8'hFF;
            14'h2F24: rddata <= 8'hFF; 14'h2F25: rddata <= 8'hFF; 14'h2F26: rddata <= 8'hFF; 14'h2F27: rddata <= 8'hFF;
            14'h2F28: rddata <= 8'hFF; 14'h2F29: rddata <= 8'hFF; 14'h2F2A: rddata <= 8'hFF; 14'h2F2B: rddata <= 8'hFF;
            14'h2F2C: rddata <= 8'hFF; 14'h2F2D: rddata <= 8'hFF; 14'h2F2E: rddata <= 8'hFF; 14'h2F2F: rddata <= 8'hFF;
            14'h2F30: rddata <= 8'hFF; 14'h2F31: rddata <= 8'hFF; 14'h2F32: rddata <= 8'hFF; 14'h2F33: rddata <= 8'hFF;
            14'h2F34: rddata <= 8'hFF; 14'h2F35: rddata <= 8'hFF; 14'h2F36: rddata <= 8'hFF; 14'h2F37: rddata <= 8'hFF;
            14'h2F38: rddata <= 8'hFF; 14'h2F39: rddata <= 8'hFF; 14'h2F3A: rddata <= 8'hFF; 14'h2F3B: rddata <= 8'hFF;
            14'h2F3C: rddata <= 8'hFF; 14'h2F3D: rddata <= 8'hFF; 14'h2F3E: rddata <= 8'hFF; 14'h2F3F: rddata <= 8'hFF;
            14'h2F40: rddata <= 8'hFF; 14'h2F41: rddata <= 8'hFF; 14'h2F42: rddata <= 8'hFF; 14'h2F43: rddata <= 8'hFF;
            14'h2F44: rddata <= 8'hFF; 14'h2F45: rddata <= 8'hFF; 14'h2F46: rddata <= 8'hFF; 14'h2F47: rddata <= 8'hFF;
            14'h2F48: rddata <= 8'hFF; 14'h2F49: rddata <= 8'hFF; 14'h2F4A: rddata <= 8'hFF; 14'h2F4B: rddata <= 8'hFF;
            14'h2F4C: rddata <= 8'hFF; 14'h2F4D: rddata <= 8'hFF; 14'h2F4E: rddata <= 8'hFF; 14'h2F4F: rddata <= 8'hFF;
            14'h2F50: rddata <= 8'hFF; 14'h2F51: rddata <= 8'hFF; 14'h2F52: rddata <= 8'hFF; 14'h2F53: rddata <= 8'hFF;
            14'h2F54: rddata <= 8'hFF; 14'h2F55: rddata <= 8'hFF; 14'h2F56: rddata <= 8'hFF; 14'h2F57: rddata <= 8'hFF;
            14'h2F58: rddata <= 8'hFF; 14'h2F59: rddata <= 8'hFF; 14'h2F5A: rddata <= 8'hFF; 14'h2F5B: rddata <= 8'hFF;
            14'h2F5C: rddata <= 8'hFF; 14'h2F5D: rddata <= 8'hFF; 14'h2F5E: rddata <= 8'hFF; 14'h2F5F: rddata <= 8'hFF;
            14'h2F60: rddata <= 8'hFF; 14'h2F61: rddata <= 8'hFF; 14'h2F62: rddata <= 8'hFF; 14'h2F63: rddata <= 8'hFF;
            14'h2F64: rddata <= 8'hFF; 14'h2F65: rddata <= 8'hFF; 14'h2F66: rddata <= 8'hFF; 14'h2F67: rddata <= 8'hFF;
            14'h2F68: rddata <= 8'hFF; 14'h2F69: rddata <= 8'hFF; 14'h2F6A: rddata <= 8'hFF; 14'h2F6B: rddata <= 8'hFF;
            14'h2F6C: rddata <= 8'hFF; 14'h2F6D: rddata <= 8'hFF; 14'h2F6E: rddata <= 8'hFF; 14'h2F6F: rddata <= 8'hFF;
            14'h2F70: rddata <= 8'hFF; 14'h2F71: rddata <= 8'hFF; 14'h2F72: rddata <= 8'hFF; 14'h2F73: rddata <= 8'hFF;
            14'h2F74: rddata <= 8'hFF; 14'h2F75: rddata <= 8'hFF; 14'h2F76: rddata <= 8'hFF; 14'h2F77: rddata <= 8'hFF;
            14'h2F78: rddata <= 8'hFF; 14'h2F79: rddata <= 8'hFF; 14'h2F7A: rddata <= 8'hFF; 14'h2F7B: rddata <= 8'hFF;
            14'h2F7C: rddata <= 8'hFF; 14'h2F7D: rddata <= 8'hFF; 14'h2F7E: rddata <= 8'hFF; 14'h2F7F: rddata <= 8'hFF;
            14'h2F80: rddata <= 8'hFF; 14'h2F81: rddata <= 8'hFF; 14'h2F82: rddata <= 8'hFF; 14'h2F83: rddata <= 8'hFF;
            14'h2F84: rddata <= 8'hFF; 14'h2F85: rddata <= 8'hFF; 14'h2F86: rddata <= 8'hFF; 14'h2F87: rddata <= 8'hFF;
            14'h2F88: rddata <= 8'hFF; 14'h2F89: rddata <= 8'hFF; 14'h2F8A: rddata <= 8'hFF; 14'h2F8B: rddata <= 8'hFF;
            14'h2F8C: rddata <= 8'hFF; 14'h2F8D: rddata <= 8'hFF; 14'h2F8E: rddata <= 8'hFF; 14'h2F8F: rddata <= 8'hFF;
            14'h2F90: rddata <= 8'hFF; 14'h2F91: rddata <= 8'hFF; 14'h2F92: rddata <= 8'hFF; 14'h2F93: rddata <= 8'hFF;
            14'h2F94: rddata <= 8'hFF; 14'h2F95: rddata <= 8'hFF; 14'h2F96: rddata <= 8'hFF; 14'h2F97: rddata <= 8'hFF;
            14'h2F98: rddata <= 8'hFF; 14'h2F99: rddata <= 8'hFF; 14'h2F9A: rddata <= 8'hFF; 14'h2F9B: rddata <= 8'hFF;
            14'h2F9C: rddata <= 8'hFF; 14'h2F9D: rddata <= 8'hFF; 14'h2F9E: rddata <= 8'hFF; 14'h2F9F: rddata <= 8'hFF;
            14'h2FA0: rddata <= 8'hFF; 14'h2FA1: rddata <= 8'hFF; 14'h2FA2: rddata <= 8'hFF; 14'h2FA3: rddata <= 8'hFF;
            14'h2FA4: rddata <= 8'hFF; 14'h2FA5: rddata <= 8'hFF; 14'h2FA6: rddata <= 8'hFF; 14'h2FA7: rddata <= 8'hFF;
            14'h2FA8: rddata <= 8'hFF; 14'h2FA9: rddata <= 8'hFF; 14'h2FAA: rddata <= 8'hFF; 14'h2FAB: rddata <= 8'hFF;
            14'h2FAC: rddata <= 8'hFF; 14'h2FAD: rddata <= 8'hFF; 14'h2FAE: rddata <= 8'hFF; 14'h2FAF: rddata <= 8'hFF;
            14'h2FB0: rddata <= 8'hFF; 14'h2FB1: rddata <= 8'hFF; 14'h2FB2: rddata <= 8'hFF; 14'h2FB3: rddata <= 8'hFF;
            14'h2FB4: rddata <= 8'hFF; 14'h2FB5: rddata <= 8'hFF; 14'h2FB6: rddata <= 8'hFF; 14'h2FB7: rddata <= 8'hFF;
            14'h2FB8: rddata <= 8'hFF; 14'h2FB9: rddata <= 8'hFF; 14'h2FBA: rddata <= 8'hFF; 14'h2FBB: rddata <= 8'hFF;
            14'h2FBC: rddata <= 8'hFF; 14'h2FBD: rddata <= 8'hFF; 14'h2FBE: rddata <= 8'hFF; 14'h2FBF: rddata <= 8'hFF;
            14'h2FC0: rddata <= 8'hFF; 14'h2FC1: rddata <= 8'hFF; 14'h2FC2: rddata <= 8'hFF; 14'h2FC3: rddata <= 8'hFF;
            14'h2FC4: rddata <= 8'hFF; 14'h2FC5: rddata <= 8'hFF; 14'h2FC6: rddata <= 8'hFF; 14'h2FC7: rddata <= 8'hFF;
            14'h2FC8: rddata <= 8'hFF; 14'h2FC9: rddata <= 8'hFF; 14'h2FCA: rddata <= 8'hFF; 14'h2FCB: rddata <= 8'hFF;
            14'h2FCC: rddata <= 8'hFF; 14'h2FCD: rddata <= 8'hFF; 14'h2FCE: rddata <= 8'hFF; 14'h2FCF: rddata <= 8'hFF;
            14'h2FD0: rddata <= 8'hFF; 14'h2FD1: rddata <= 8'hFF; 14'h2FD2: rddata <= 8'hFF; 14'h2FD3: rddata <= 8'hFF;
            14'h2FD4: rddata <= 8'hFF; 14'h2FD5: rddata <= 8'hFF; 14'h2FD6: rddata <= 8'hFF; 14'h2FD7: rddata <= 8'hFF;
            14'h2FD8: rddata <= 8'hFF; 14'h2FD9: rddata <= 8'hFF; 14'h2FDA: rddata <= 8'hFF; 14'h2FDB: rddata <= 8'hFF;
            14'h2FDC: rddata <= 8'hFF; 14'h2FDD: rddata <= 8'hFF; 14'h2FDE: rddata <= 8'hFF; 14'h2FDF: rddata <= 8'hFF;
            14'h2FE0: rddata <= 8'hFF; 14'h2FE1: rddata <= 8'hFF; 14'h2FE2: rddata <= 8'hFF; 14'h2FE3: rddata <= 8'hFF;
            14'h2FE4: rddata <= 8'hFF; 14'h2FE5: rddata <= 8'hFF; 14'h2FE6: rddata <= 8'hFF; 14'h2FE7: rddata <= 8'hFF;
            14'h2FE8: rddata <= 8'hFF; 14'h2FE9: rddata <= 8'hFF; 14'h2FEA: rddata <= 8'hFF; 14'h2FEB: rddata <= 8'hFF;
            14'h2FEC: rddata <= 8'hFF; 14'h2FED: rddata <= 8'hFF; 14'h2FEE: rddata <= 8'hFF; 14'h2FEF: rddata <= 8'hFF;
            14'h2FF0: rddata <= 8'hFF; 14'h2FF1: rddata <= 8'hFF; 14'h2FF2: rddata <= 8'hFF; 14'h2FF3: rddata <= 8'hFF;
            14'h2FF4: rddata <= 8'hFF; 14'h2FF5: rddata <= 8'hFF; 14'h2FF6: rddata <= 8'hFF; 14'h2FF7: rddata <= 8'hFF;
            14'h2FF8: rddata <= 8'hFF; 14'h2FF9: rddata <= 8'hFF; 14'h2FFA: rddata <= 8'hFF; 14'h2FFB: rddata <= 8'hFF;
            14'h2FFC: rddata <= 8'hFF; 14'h2FFD: rddata <= 8'hFF; 14'h2FFE: rddata <= 8'hFF; 14'h2FFF: rddata <= 8'hFF;
            14'h3000: rddata <= 8'h3C; 14'h3001: rddata <= 8'h20; 14'h3002: rddata <= 8'h20; 14'h3003: rddata <= 8'h78;
            14'h3004: rddata <= 8'h20; 14'h3005: rddata <= 8'h60; 14'h3006: rddata <= 8'hAC; 14'h3007: rddata <= 8'h00;
            14'h3008: rddata <= 8'h44; 14'h3009: rddata <= 8'h48; 14'h300A: rddata <= 8'h50; 14'h300B: rddata <= 8'h2C;
            14'h300C: rddata <= 8'h44; 14'h300D: rddata <= 8'h08; 14'h300E: rddata <= 8'h1C; 14'h300F: rddata <= 8'h00;
            14'h3010: rddata <= 8'h44; 14'h3011: rddata <= 8'h48; 14'h3012: rddata <= 8'h50; 14'h3013: rddata <= 8'h2C;
            14'h3014: rddata <= 8'h54; 14'h3015: rddata <= 8'h1C; 14'h3016: rddata <= 8'h04; 14'h3017: rddata <= 8'h00;
            14'h3018: rddata <= 8'h64; 14'h3019: rddata <= 8'h28; 14'h301A: rddata <= 8'h50; 14'h301B: rddata <= 8'h2C;
            14'h301C: rddata <= 8'h54; 14'h301D: rddata <= 8'h1C; 14'h301E: rddata <= 8'h04; 14'h301F: rddata <= 8'h00;
            14'h3020: rddata <= 8'h00; 14'h3021: rddata <= 8'h10; 14'h3022: rddata <= 8'h00; 14'h3023: rddata <= 8'h7C;
            14'h3024: rddata <= 8'h00; 14'h3025: rddata <= 8'h10; 14'h3026: rddata <= 8'h00; 14'h3027: rddata <= 8'h00;
            14'h3028: rddata <= 8'h3C; 14'h3029: rddata <= 8'h42; 14'h302A: rddata <= 8'h99; 14'h302B: rddata <= 8'hA1;
            14'h302C: rddata <= 8'hA1; 14'h302D: rddata <= 8'h99; 14'h302E: rddata <= 8'h42; 14'h302F: rddata <= 8'h3C;
            14'h3030: rddata <= 8'h00; 14'h3031: rddata <= 8'h04; 14'h3032: rddata <= 8'h02; 14'h3033: rddata <= 8'hFF;
            14'h3034: rddata <= 8'hFF; 14'h3035: rddata <= 8'h02; 14'h3036: rddata <= 8'h04; 14'h3037: rddata <= 8'h00;
            14'h3038: rddata <= 8'h00; 14'h3039: rddata <= 8'h20; 14'h303A: rddata <= 8'h40; 14'h303B: rddata <= 8'hFF;
            14'h303C: rddata <= 8'hFF; 14'h303D: rddata <= 8'h40; 14'h303E: rddata <= 8'h20; 14'h303F: rddata <= 8'h00;
            14'h3040: rddata <= 8'h18; 14'h3041: rddata <= 8'h3C; 14'h3042: rddata <= 8'h5A; 14'h3043: rddata <= 8'h18;
            14'h3044: rddata <= 8'h18; 14'h3045: rddata <= 8'h18; 14'h3046: rddata <= 8'h18; 14'h3047: rddata <= 8'h18;
            14'h3048: rddata <= 8'h18; 14'h3049: rddata <= 8'h18; 14'h304A: rddata <= 8'h18; 14'h304B: rddata <= 8'h18;
            14'h304C: rddata <= 8'h18; 14'h304D: rddata <= 8'h5A; 14'h304E: rddata <= 8'h3C; 14'h304F: rddata <= 8'h18;
            14'h3050: rddata <= 8'h0F; 14'h3051: rddata <= 8'h07; 14'h3052: rddata <= 8'h0F; 14'h3053: rddata <= 8'h1D;
            14'h3054: rddata <= 8'h38; 14'h3055: rddata <= 8'h70; 14'h3056: rddata <= 8'h20; 14'h3057: rddata <= 8'h00;
            14'h3058: rddata <= 8'h00; 14'h3059: rddata <= 8'h04; 14'h305A: rddata <= 8'h0E; 14'h305B: rddata <= 8'h1C;
            14'h305C: rddata <= 8'hB8; 14'h305D: rddata <= 8'hF0; 14'h305E: rddata <= 8'hE0; 14'h305F: rddata <= 8'hF0;
            14'h3060: rddata <= 8'h00; 14'h3061: rddata <= 8'h20; 14'h3062: rddata <= 8'h70; 14'h3063: rddata <= 8'h38;
            14'h3064: rddata <= 8'h1D; 14'h3065: rddata <= 8'h0F; 14'h3066: rddata <= 8'h07; 14'h3067: rddata <= 8'h0F;
            14'h3068: rddata <= 8'hF0; 14'h3069: rddata <= 8'hE0; 14'h306A: rddata <= 8'hF0; 14'h306B: rddata <= 8'hB8;
            14'h306C: rddata <= 8'h1C; 14'h306D: rddata <= 8'h0E; 14'h306E: rddata <= 8'h04; 14'h306F: rddata <= 8'h00;
            14'h3070: rddata <= 8'h00; 14'h3071: rddata <= 8'h3C; 14'h3072: rddata <= 8'h3C; 14'h3073: rddata <= 8'h00;
            14'h3074: rddata <= 8'h7E; 14'h3075: rddata <= 8'hFF; 14'h3076: rddata <= 8'hFF; 14'h3077: rddata <= 8'hFF;
            14'h3078: rddata <= 8'hFC; 14'h3079: rddata <= 8'hFC; 14'h307A: rddata <= 8'h3C; 14'h307B: rddata <= 8'h30;
            14'h307C: rddata <= 8'h30; 14'h307D: rddata <= 8'h30; 14'h307E: rddata <= 8'h30; 14'h307F: rddata <= 8'h30;
            14'h3080: rddata <= 8'hFF; 14'h3081: rddata <= 8'h3C; 14'h3082: rddata <= 8'h3C; 14'h3083: rddata <= 8'h3C;
            14'h3084: rddata <= 8'h3C; 14'h3085: rddata <= 8'h00; 14'h3086: rddata <= 8'h00; 14'h3087: rddata <= 8'h00;
            14'h3088: rddata <= 8'h3F; 14'h3089: rddata <= 8'h3F; 14'h308A: rddata <= 8'h3C; 14'h308B: rddata <= 8'h0C;
            14'h308C: rddata <= 8'h0C; 14'h308D: rddata <= 8'h0C; 14'h308E: rddata <= 8'h0C; 14'h308F: rddata <= 8'h0C;
            14'h3090: rddata <= 8'h3C; 14'h3091: rddata <= 8'h3C; 14'h3092: rddata <= 8'h3C; 14'h3093: rddata <= 8'h3C;
            14'h3094: rddata <= 8'h3C; 14'h3095: rddata <= 8'h3C; 14'h3096: rddata <= 8'h3C; 14'h3097: rddata <= 8'h3C;
            14'h3098: rddata <= 8'h00; 14'h3099: rddata <= 8'h3C; 14'h309A: rddata <= 8'h3C; 14'h309B: rddata <= 8'h00;
            14'h309C: rddata <= 8'h7E; 14'h309D: rddata <= 8'hFF; 14'h309E: rddata <= 8'hBD; 14'h309F: rddata <= 8'hDB;
            14'h30A0: rddata <= 8'h7E; 14'h30A1: rddata <= 8'h3C; 14'h30A2: rddata <= 8'h66; 14'h30A3: rddata <= 8'h66;
            14'h30A4: rddata <= 8'hE7; 14'h30A5: rddata <= 8'hC3; 14'h30A6: rddata <= 8'hC3; 14'h30A7: rddata <= 8'hC3;
            14'h30A8: rddata <= 8'h00; 14'h30A9: rddata <= 8'h38; 14'h30AA: rddata <= 8'h3C; 14'h30AB: rddata <= 8'h00;
            14'h30AC: rddata <= 8'h38; 14'h30AD: rddata <= 8'h78; 14'h30AE: rddata <= 8'h7C; 14'h30AF: rddata <= 8'h7F;
            14'h30B0: rddata <= 8'h7C; 14'h30B1: rddata <= 8'h3E; 14'h30B2: rddata <= 8'h1B; 14'h30B3: rddata <= 8'h1E;
            14'h30B4: rddata <= 8'h1C; 14'h30B5: rddata <= 8'h18; 14'h30B6: rddata <= 8'h38; 14'h30B7: rddata <= 8'h38;
            14'h30B8: rddata <= 8'h00; 14'h30B9: rddata <= 8'h38; 14'h30BA: rddata <= 8'h3C; 14'h30BB: rddata <= 8'h00;
            14'h30BC: rddata <= 8'h39; 14'h30BD: rddata <= 8'h79; 14'h30BE: rddata <= 8'hDF; 14'h30BF: rddata <= 8'hDC;
            14'h30C0: rddata <= 8'h7C; 14'h30C1: rddata <= 8'h3F; 14'h30C2: rddata <= 8'h1F; 14'h30C3: rddata <= 8'h3B;
            14'h30C4: rddata <= 8'hF3; 14'h30C5: rddata <= 8'hC3; 14'h30C6: rddata <= 8'h80; 14'h30C7: rddata <= 8'h00;
            14'h30C8: rddata <= 8'h18; 14'h30C9: rddata <= 8'h3C; 14'h30CA: rddata <= 8'h66; 14'h30CB: rddata <= 8'h24;
            14'h30CC: rddata <= 8'hE7; 14'h30CD: rddata <= 8'hBD; 14'h30CE: rddata <= 8'h99; 14'h30CF: rddata <= 8'hDB;
            14'h30D0: rddata <= 8'h00; 14'h30D1: rddata <= 8'h00; 14'h30D2: rddata <= 8'h00; 14'h30D3: rddata <= 8'h00;
            14'h30D4: rddata <= 8'h0F; 14'h30D5: rddata <= 8'h0F; 14'h30D6: rddata <= 8'h0F; 14'h30D7: rddata <= 8'h0F;
            14'h30D8: rddata <= 8'h0F; 14'h30D9: rddata <= 8'h0F; 14'h30DA: rddata <= 8'h0F; 14'h30DB: rddata <= 8'h0F;
            14'h30DC: rddata <= 8'h00; 14'h30DD: rddata <= 8'h00; 14'h30DE: rddata <= 8'h00; 14'h30DF: rddata <= 8'h00;
            14'h30E0: rddata <= 8'h00; 14'h30E1: rddata <= 8'h00; 14'h30E2: rddata <= 8'h00; 14'h30E3: rddata <= 8'h00;
            14'h30E4: rddata <= 8'hF0; 14'h30E5: rddata <= 8'hF0; 14'h30E6: rddata <= 8'hF0; 14'h30E7: rddata <= 8'hF0;
            14'h30E8: rddata <= 8'hF0; 14'h30E9: rddata <= 8'hF0; 14'h30EA: rddata <= 8'hF0; 14'h30EB: rddata <= 8'hF0;
            14'h30EC: rddata <= 8'h00; 14'h30ED: rddata <= 8'h00; 14'h30EE: rddata <= 8'h00; 14'h30EF: rddata <= 8'h00;
            14'h30F0: rddata <= 8'hF0; 14'h30F1: rddata <= 8'hF0; 14'h30F2: rddata <= 8'hF0; 14'h30F3: rddata <= 8'hF0;
            14'h30F4: rddata <= 8'h0F; 14'h30F5: rddata <= 8'h0F; 14'h30F6: rddata <= 8'h0F; 14'h30F7: rddata <= 8'h0F;
            14'h30F8: rddata <= 8'h00; 14'h30F9: rddata <= 8'h00; 14'h30FA: rddata <= 8'h00; 14'h30FB: rddata <= 8'h00;
            14'h30FC: rddata <= 8'hFF; 14'h30FD: rddata <= 8'hFF; 14'h30FE: rddata <= 8'hFF; 14'h30FF: rddata <= 8'hFF;
            14'h3100: rddata <= 8'h00; 14'h3101: rddata <= 8'h00; 14'h3102: rddata <= 8'h00; 14'h3103: rddata <= 8'h00;
            14'h3104: rddata <= 8'h00; 14'h3105: rddata <= 8'h00; 14'h3106: rddata <= 8'h00; 14'h3107: rddata <= 8'h00;
            14'h3108: rddata <= 8'h10; 14'h3109: rddata <= 8'h10; 14'h310A: rddata <= 8'h10; 14'h310B: rddata <= 8'h10;
            14'h310C: rddata <= 8'h10; 14'h310D: rddata <= 8'h00; 14'h310E: rddata <= 8'h10; 14'h310F: rddata <= 8'h00;
            14'h3110: rddata <= 8'h28; 14'h3111: rddata <= 8'h28; 14'h3112: rddata <= 8'h28; 14'h3113: rddata <= 8'h00;
            14'h3114: rddata <= 8'h00; 14'h3115: rddata <= 8'h00; 14'h3116: rddata <= 8'h00; 14'h3117: rddata <= 8'h00;
            14'h3118: rddata <= 8'h28; 14'h3119: rddata <= 8'h28; 14'h311A: rddata <= 8'h7C; 14'h311B: rddata <= 8'h28;
            14'h311C: rddata <= 8'h7C; 14'h311D: rddata <= 8'h28; 14'h311E: rddata <= 8'h28; 14'h311F: rddata <= 8'h00;
            14'h3120: rddata <= 8'h10; 14'h3121: rddata <= 8'h3C; 14'h3122: rddata <= 8'h50; 14'h3123: rddata <= 8'h38;
            14'h3124: rddata <= 8'h14; 14'h3125: rddata <= 8'h78; 14'h3126: rddata <= 8'h10; 14'h3127: rddata <= 8'h00;
            14'h3128: rddata <= 8'h60; 14'h3129: rddata <= 8'h64; 14'h312A: rddata <= 8'h08; 14'h312B: rddata <= 8'h10;
            14'h312C: rddata <= 8'h20; 14'h312D: rddata <= 8'h4C; 14'h312E: rddata <= 8'h0C; 14'h312F: rddata <= 8'h00;
            14'h3130: rddata <= 8'h20; 14'h3131: rddata <= 8'h50; 14'h3132: rddata <= 8'h50; 14'h3133: rddata <= 8'h20;
            14'h3134: rddata <= 8'h54; 14'h3135: rddata <= 8'h48; 14'h3136: rddata <= 8'h34; 14'h3137: rddata <= 8'h00;
            14'h3138: rddata <= 8'h08; 14'h3139: rddata <= 8'h08; 14'h313A: rddata <= 8'h10; 14'h313B: rddata <= 8'h00;
            14'h313C: rddata <= 8'h00; 14'h313D: rddata <= 8'h00; 14'h313E: rddata <= 8'h00; 14'h313F: rddata <= 8'h00;
            14'h3140: rddata <= 8'h10; 14'h3141: rddata <= 8'h20; 14'h3142: rddata <= 8'h40; 14'h3143: rddata <= 8'h40;
            14'h3144: rddata <= 8'h40; 14'h3145: rddata <= 8'h20; 14'h3146: rddata <= 8'h10; 14'h3147: rddata <= 8'h00;
            14'h3148: rddata <= 8'h10; 14'h3149: rddata <= 8'h08; 14'h314A: rddata <= 8'h04; 14'h314B: rddata <= 8'h04;
            14'h314C: rddata <= 8'h04; 14'h314D: rddata <= 8'h08; 14'h314E: rddata <= 8'h10; 14'h314F: rddata <= 8'h00;
            14'h3150: rddata <= 8'h10; 14'h3151: rddata <= 8'h54; 14'h3152: rddata <= 8'h38; 14'h3153: rddata <= 8'h10;
            14'h3154: rddata <= 8'h38; 14'h3155: rddata <= 8'h54; 14'h3156: rddata <= 8'h10; 14'h3157: rddata <= 8'h00;
            14'h3158: rddata <= 8'h00; 14'h3159: rddata <= 8'h10; 14'h315A: rddata <= 8'h10; 14'h315B: rddata <= 8'h7C;
            14'h315C: rddata <= 8'h10; 14'h315D: rddata <= 8'h10; 14'h315E: rddata <= 8'h00; 14'h315F: rddata <= 8'h00;
            14'h3160: rddata <= 8'h00; 14'h3161: rddata <= 8'h00; 14'h3162: rddata <= 8'h00; 14'h3163: rddata <= 8'h00;
            14'h3164: rddata <= 8'h10; 14'h3165: rddata <= 8'h10; 14'h3166: rddata <= 8'h20; 14'h3167: rddata <= 8'h00;
            14'h3168: rddata <= 8'h00; 14'h3169: rddata <= 8'h00; 14'h316A: rddata <= 8'h00; 14'h316B: rddata <= 8'h7C;
            14'h316C: rddata <= 8'h00; 14'h316D: rddata <= 8'h00; 14'h316E: rddata <= 8'h00; 14'h316F: rddata <= 8'h00;
            14'h3170: rddata <= 8'h00; 14'h3171: rddata <= 8'h00; 14'h3172: rddata <= 8'h00; 14'h3173: rddata <= 8'h00;
            14'h3174: rddata <= 8'h00; 14'h3175: rddata <= 8'h00; 14'h3176: rddata <= 8'h10; 14'h3177: rddata <= 8'h00;
            14'h3178: rddata <= 8'h00; 14'h3179: rddata <= 8'h04; 14'h317A: rddata <= 8'h08; 14'h317B: rddata <= 8'h10;
            14'h317C: rddata <= 8'h20; 14'h317D: rddata <= 8'h40; 14'h317E: rddata <= 8'h00; 14'h317F: rddata <= 8'h00;
            14'h3180: rddata <= 8'h38; 14'h3181: rddata <= 8'h44; 14'h3182: rddata <= 8'h4C; 14'h3183: rddata <= 8'h54;
            14'h3184: rddata <= 8'h64; 14'h3185: rddata <= 8'h44; 14'h3186: rddata <= 8'h38; 14'h3187: rddata <= 8'h00;
            14'h3188: rddata <= 8'h10; 14'h3189: rddata <= 8'h30; 14'h318A: rddata <= 8'h10; 14'h318B: rddata <= 8'h10;
            14'h318C: rddata <= 8'h10; 14'h318D: rddata <= 8'h10; 14'h318E: rddata <= 8'h38; 14'h318F: rddata <= 8'h00;
            14'h3190: rddata <= 8'h38; 14'h3191: rddata <= 8'h44; 14'h3192: rddata <= 8'h04; 14'h3193: rddata <= 8'h18;
            14'h3194: rddata <= 8'h20; 14'h3195: rddata <= 8'h40; 14'h3196: rddata <= 8'h7C; 14'h3197: rddata <= 8'h00;
            14'h3198: rddata <= 8'h7C; 14'h3199: rddata <= 8'h04; 14'h319A: rddata <= 8'h08; 14'h319B: rddata <= 8'h18;
            14'h319C: rddata <= 8'h04; 14'h319D: rddata <= 8'h44; 14'h319E: rddata <= 8'h38; 14'h319F: rddata <= 8'h00;
            14'h31A0: rddata <= 8'h08; 14'h31A1: rddata <= 8'h18; 14'h31A2: rddata <= 8'h28; 14'h31A3: rddata <= 8'h48;
            14'h31A4: rddata <= 8'h7C; 14'h31A5: rddata <= 8'h08; 14'h31A6: rddata <= 8'h08; 14'h31A7: rddata <= 8'h00;
            14'h31A8: rddata <= 8'h7C; 14'h31A9: rddata <= 8'h40; 14'h31AA: rddata <= 8'h78; 14'h31AB: rddata <= 8'h04;
            14'h31AC: rddata <= 8'h04; 14'h31AD: rddata <= 8'h44; 14'h31AE: rddata <= 8'h38; 14'h31AF: rddata <= 8'h00;
            14'h31B0: rddata <= 8'h1C; 14'h31B1: rddata <= 8'h20; 14'h31B2: rddata <= 8'h40; 14'h31B3: rddata <= 8'h78;
            14'h31B4: rddata <= 8'h44; 14'h31B5: rddata <= 8'h44; 14'h31B6: rddata <= 8'h38; 14'h31B7: rddata <= 8'h00;
            14'h31B8: rddata <= 8'h7C; 14'h31B9: rddata <= 8'h04; 14'h31BA: rddata <= 8'h08; 14'h31BB: rddata <= 8'h10;
            14'h31BC: rddata <= 8'h20; 14'h31BD: rddata <= 8'h20; 14'h31BE: rddata <= 8'h20; 14'h31BF: rddata <= 8'h00;
            14'h31C0: rddata <= 8'h38; 14'h31C1: rddata <= 8'h44; 14'h31C2: rddata <= 8'h44; 14'h31C3: rddata <= 8'h38;
            14'h31C4: rddata <= 8'h44; 14'h31C5: rddata <= 8'h44; 14'h31C6: rddata <= 8'h38; 14'h31C7: rddata <= 8'h00;
            14'h31C8: rddata <= 8'h38; 14'h31C9: rddata <= 8'h44; 14'h31CA: rddata <= 8'h44; 14'h31CB: rddata <= 8'h3C;
            14'h31CC: rddata <= 8'h04; 14'h31CD: rddata <= 8'h08; 14'h31CE: rddata <= 8'h70; 14'h31CF: rddata <= 8'h00;
            14'h31D0: rddata <= 8'h00; 14'h31D1: rddata <= 8'h00; 14'h31D2: rddata <= 8'h10; 14'h31D3: rddata <= 8'h00;
            14'h31D4: rddata <= 8'h10; 14'h31D5: rddata <= 8'h00; 14'h31D6: rddata <= 8'h00; 14'h31D7: rddata <= 8'h00;
            14'h31D8: rddata <= 8'h00; 14'h31D9: rddata <= 8'h00; 14'h31DA: rddata <= 8'h10; 14'h31DB: rddata <= 8'h00;
            14'h31DC: rddata <= 8'h10; 14'h31DD: rddata <= 8'h10; 14'h31DE: rddata <= 8'h20; 14'h31DF: rddata <= 8'h00;
            14'h31E0: rddata <= 8'h08; 14'h31E1: rddata <= 8'h10; 14'h31E2: rddata <= 8'h20; 14'h31E3: rddata <= 8'h40;
            14'h31E4: rddata <= 8'h20; 14'h31E5: rddata <= 8'h10; 14'h31E6: rddata <= 8'h08; 14'h31E7: rddata <= 8'h00;
            14'h31E8: rddata <= 8'h00; 14'h31E9: rddata <= 8'h00; 14'h31EA: rddata <= 8'h7C; 14'h31EB: rddata <= 8'h00;
            14'h31EC: rddata <= 8'h7C; 14'h31ED: rddata <= 8'h00; 14'h31EE: rddata <= 8'h00; 14'h31EF: rddata <= 8'h00;
            14'h31F0: rddata <= 8'h20; 14'h31F1: rddata <= 8'h10; 14'h31F2: rddata <= 8'h08; 14'h31F3: rddata <= 8'h04;
            14'h31F4: rddata <= 8'h08; 14'h31F5: rddata <= 8'h10; 14'h31F6: rddata <= 8'h20; 14'h31F7: rddata <= 8'h00;
            14'h31F8: rddata <= 8'h38; 14'h31F9: rddata <= 8'h44; 14'h31FA: rddata <= 8'h08; 14'h31FB: rddata <= 8'h10;
            14'h31FC: rddata <= 8'h10; 14'h31FD: rddata <= 8'h00; 14'h31FE: rddata <= 8'h10; 14'h31FF: rddata <= 8'h00;
            14'h3200: rddata <= 8'h38; 14'h3201: rddata <= 8'h44; 14'h3202: rddata <= 8'h54; 14'h3203: rddata <= 8'h5C;
            14'h3204: rddata <= 8'h58; 14'h3205: rddata <= 8'h40; 14'h3206: rddata <= 8'h3C; 14'h3207: rddata <= 8'h00;
            14'h3208: rddata <= 8'h10; 14'h3209: rddata <= 8'h28; 14'h320A: rddata <= 8'h44; 14'h320B: rddata <= 8'h44;
            14'h320C: rddata <= 8'h7C; 14'h320D: rddata <= 8'h44; 14'h320E: rddata <= 8'h44; 14'h320F: rddata <= 8'h00;
            14'h3210: rddata <= 8'h78; 14'h3211: rddata <= 8'h44; 14'h3212: rddata <= 8'h44; 14'h3213: rddata <= 8'h78;
            14'h3214: rddata <= 8'h44; 14'h3215: rddata <= 8'h44; 14'h3216: rddata <= 8'h78; 14'h3217: rddata <= 8'h00;
            14'h3218: rddata <= 8'h38; 14'h3219: rddata <= 8'h44; 14'h321A: rddata <= 8'h40; 14'h321B: rddata <= 8'h40;
            14'h321C: rddata <= 8'h40; 14'h321D: rddata <= 8'h44; 14'h321E: rddata <= 8'h38; 14'h321F: rddata <= 8'h00;
            14'h3220: rddata <= 8'h78; 14'h3221: rddata <= 8'h44; 14'h3222: rddata <= 8'h44; 14'h3223: rddata <= 8'h44;
            14'h3224: rddata <= 8'h44; 14'h3225: rddata <= 8'h44; 14'h3226: rddata <= 8'h78; 14'h3227: rddata <= 8'h00;
            14'h3228: rddata <= 8'h7C; 14'h3229: rddata <= 8'h40; 14'h322A: rddata <= 8'h40; 14'h322B: rddata <= 8'h78;
            14'h322C: rddata <= 8'h40; 14'h322D: rddata <= 8'h40; 14'h322E: rddata <= 8'h7C; 14'h322F: rddata <= 8'h00;
            14'h3230: rddata <= 8'h7C; 14'h3231: rddata <= 8'h40; 14'h3232: rddata <= 8'h40; 14'h3233: rddata <= 8'h78;
            14'h3234: rddata <= 8'h40; 14'h3235: rddata <= 8'h40; 14'h3236: rddata <= 8'h40; 14'h3237: rddata <= 8'h00;
            14'h3238: rddata <= 8'h3C; 14'h3239: rddata <= 8'h40; 14'h323A: rddata <= 8'h40; 14'h323B: rddata <= 8'h40;
            14'h323C: rddata <= 8'h4C; 14'h323D: rddata <= 8'h44; 14'h323E: rddata <= 8'h3C; 14'h323F: rddata <= 8'h00;
            14'h3240: rddata <= 8'h44; 14'h3241: rddata <= 8'h44; 14'h3242: rddata <= 8'h44; 14'h3243: rddata <= 8'h7C;
            14'h3244: rddata <= 8'h44; 14'h3245: rddata <= 8'h44; 14'h3246: rddata <= 8'h44; 14'h3247: rddata <= 8'h00;
            14'h3248: rddata <= 8'h38; 14'h3249: rddata <= 8'h10; 14'h324A: rddata <= 8'h10; 14'h324B: rddata <= 8'h10;
            14'h324C: rddata <= 8'h10; 14'h324D: rddata <= 8'h10; 14'h324E: rddata <= 8'h38; 14'h324F: rddata <= 8'h00;
            14'h3250: rddata <= 8'h04; 14'h3251: rddata <= 8'h04; 14'h3252: rddata <= 8'h04; 14'h3253: rddata <= 8'h04;
            14'h3254: rddata <= 8'h04; 14'h3255: rddata <= 8'h44; 14'h3256: rddata <= 8'h38; 14'h3257: rddata <= 8'h00;
            14'h3258: rddata <= 8'h44; 14'h3259: rddata <= 8'h48; 14'h325A: rddata <= 8'h50; 14'h325B: rddata <= 8'h60;
            14'h325C: rddata <= 8'h50; 14'h325D: rddata <= 8'h48; 14'h325E: rddata <= 8'h44; 14'h325F: rddata <= 8'h00;
            14'h3260: rddata <= 8'h40; 14'h3261: rddata <= 8'h40; 14'h3262: rddata <= 8'h40; 14'h3263: rddata <= 8'h40;
            14'h3264: rddata <= 8'h40; 14'h3265: rddata <= 8'h40; 14'h3266: rddata <= 8'h7C; 14'h3267: rddata <= 8'h00;
            14'h3268: rddata <= 8'h44; 14'h3269: rddata <= 8'h6C; 14'h326A: rddata <= 8'h54; 14'h326B: rddata <= 8'h54;
            14'h326C: rddata <= 8'h44; 14'h326D: rddata <= 8'h44; 14'h326E: rddata <= 8'h44; 14'h326F: rddata <= 8'h00;
            14'h3270: rddata <= 8'h44; 14'h3271: rddata <= 8'h44; 14'h3272: rddata <= 8'h64; 14'h3273: rddata <= 8'h54;
            14'h3274: rddata <= 8'h4C; 14'h3275: rddata <= 8'h44; 14'h3276: rddata <= 8'h44; 14'h3277: rddata <= 8'h00;
            14'h3278: rddata <= 8'h38; 14'h3279: rddata <= 8'h44; 14'h327A: rddata <= 8'h44; 14'h327B: rddata <= 8'h44;
            14'h327C: rddata <= 8'h44; 14'h327D: rddata <= 8'h44; 14'h327E: rddata <= 8'h38; 14'h327F: rddata <= 8'h00;
            14'h3280: rddata <= 8'h78; 14'h3281: rddata <= 8'h44; 14'h3282: rddata <= 8'h44; 14'h3283: rddata <= 8'h78;
            14'h3284: rddata <= 8'h40; 14'h3285: rddata <= 8'h40; 14'h3286: rddata <= 8'h40; 14'h3287: rddata <= 8'h00;
            14'h3288: rddata <= 8'h38; 14'h3289: rddata <= 8'h44; 14'h328A: rddata <= 8'h44; 14'h328B: rddata <= 8'h44;
            14'h328C: rddata <= 8'h54; 14'h328D: rddata <= 8'h48; 14'h328E: rddata <= 8'h34; 14'h328F: rddata <= 8'h00;
            14'h3290: rddata <= 8'h78; 14'h3291: rddata <= 8'h44; 14'h3292: rddata <= 8'h44; 14'h3293: rddata <= 8'h78;
            14'h3294: rddata <= 8'h50; 14'h3295: rddata <= 8'h48; 14'h3296: rddata <= 8'h44; 14'h3297: rddata <= 8'h00;
            14'h3298: rddata <= 8'h38; 14'h3299: rddata <= 8'h44; 14'h329A: rddata <= 8'h40; 14'h329B: rddata <= 8'h38;
            14'h329C: rddata <= 8'h04; 14'h329D: rddata <= 8'h44; 14'h329E: rddata <= 8'h38; 14'h329F: rddata <= 8'h00;
            14'h32A0: rddata <= 8'h7C; 14'h32A1: rddata <= 8'h10; 14'h32A2: rddata <= 8'h10; 14'h32A3: rddata <= 8'h10;
            14'h32A4: rddata <= 8'h10; 14'h32A5: rddata <= 8'h10; 14'h32A6: rddata <= 8'h10; 14'h32A7: rddata <= 8'h00;
            14'h32A8: rddata <= 8'h44; 14'h32A9: rddata <= 8'h44; 14'h32AA: rddata <= 8'h44; 14'h32AB: rddata <= 8'h44;
            14'h32AC: rddata <= 8'h44; 14'h32AD: rddata <= 8'h44; 14'h32AE: rddata <= 8'h38; 14'h32AF: rddata <= 8'h00;
            14'h32B0: rddata <= 8'h44; 14'h32B1: rddata <= 8'h44; 14'h32B2: rddata <= 8'h44; 14'h32B3: rddata <= 8'h44;
            14'h32B4: rddata <= 8'h44; 14'h32B5: rddata <= 8'h28; 14'h32B6: rddata <= 8'h10; 14'h32B7: rddata <= 8'h00;
            14'h32B8: rddata <= 8'h44; 14'h32B9: rddata <= 8'h44; 14'h32BA: rddata <= 8'h44; 14'h32BB: rddata <= 8'h54;
            14'h32BC: rddata <= 8'h54; 14'h32BD: rddata <= 8'h6C; 14'h32BE: rddata <= 8'h44; 14'h32BF: rddata <= 8'h00;
            14'h32C0: rddata <= 8'h44; 14'h32C1: rddata <= 8'h44; 14'h32C2: rddata <= 8'h28; 14'h32C3: rddata <= 8'h10;
            14'h32C4: rddata <= 8'h28; 14'h32C5: rddata <= 8'h44; 14'h32C6: rddata <= 8'h44; 14'h32C7: rddata <= 8'h00;
            14'h32C8: rddata <= 8'h44; 14'h32C9: rddata <= 8'h44; 14'h32CA: rddata <= 8'h28; 14'h32CB: rddata <= 8'h10;
            14'h32CC: rddata <= 8'h10; 14'h32CD: rddata <= 8'h10; 14'h32CE: rddata <= 8'h10; 14'h32CF: rddata <= 8'h00;
            14'h32D0: rddata <= 8'h7C; 14'h32D1: rddata <= 8'h04; 14'h32D2: rddata <= 8'h08; 14'h32D3: rddata <= 8'h10;
            14'h32D4: rddata <= 8'h20; 14'h32D5: rddata <= 8'h40; 14'h32D6: rddata <= 8'h7C; 14'h32D7: rddata <= 8'h00;
            14'h32D8: rddata <= 8'h7C; 14'h32D9: rddata <= 8'h60; 14'h32DA: rddata <= 8'h60; 14'h32DB: rddata <= 8'h60;
            14'h32DC: rddata <= 8'h60; 14'h32DD: rddata <= 8'h60; 14'h32DE: rddata <= 8'h7C; 14'h32DF: rddata <= 8'h00;
            14'h32E0: rddata <= 8'h00; 14'h32E1: rddata <= 8'h40; 14'h32E2: rddata <= 8'h20; 14'h32E3: rddata <= 8'h10;
            14'h32E4: rddata <= 8'h08; 14'h32E5: rddata <= 8'h04; 14'h32E6: rddata <= 8'h00; 14'h32E7: rddata <= 8'h00;
            14'h32E8: rddata <= 8'h7C; 14'h32E9: rddata <= 8'h0C; 14'h32EA: rddata <= 8'h0C; 14'h32EB: rddata <= 8'h0C;
            14'h32EC: rddata <= 8'h0C; 14'h32ED: rddata <= 8'h0C; 14'h32EE: rddata <= 8'h7C; 14'h32EF: rddata <= 8'h00;
            14'h32F0: rddata <= 8'h00; 14'h32F1: rddata <= 8'h00; 14'h32F2: rddata <= 8'h10; 14'h32F3: rddata <= 8'h28;
            14'h32F4: rddata <= 8'h44; 14'h32F5: rddata <= 8'h00; 14'h32F6: rddata <= 8'h00; 14'h32F7: rddata <= 8'h00;
            14'h32F8: rddata <= 8'h00; 14'h32F9: rddata <= 8'h00; 14'h32FA: rddata <= 8'h00; 14'h32FB: rddata <= 8'h00;
            14'h32FC: rddata <= 8'h00; 14'h32FD: rddata <= 8'h00; 14'h32FE: rddata <= 8'h7C; 14'h32FF: rddata <= 8'h00;
            14'h3300: rddata <= 8'h20; 14'h3301: rddata <= 8'h20; 14'h3302: rddata <= 8'h10; 14'h3303: rddata <= 8'h00;
            14'h3304: rddata <= 8'h00; 14'h3305: rddata <= 8'h00; 14'h3306: rddata <= 8'h00; 14'h3307: rddata <= 8'h00;
            14'h3308: rddata <= 8'h00; 14'h3309: rddata <= 8'h00; 14'h330A: rddata <= 8'h34; 14'h330B: rddata <= 8'h4C;
            14'h330C: rddata <= 8'h44; 14'h330D: rddata <= 8'h4C; 14'h330E: rddata <= 8'h34; 14'h330F: rddata <= 8'h00;
            14'h3310: rddata <= 8'h40; 14'h3311: rddata <= 8'h40; 14'h3312: rddata <= 8'h58; 14'h3313: rddata <= 8'h64;
            14'h3314: rddata <= 8'h44; 14'h3315: rddata <= 8'h64; 14'h3316: rddata <= 8'h58; 14'h3317: rddata <= 8'h00;
            14'h3318: rddata <= 8'h00; 14'h3319: rddata <= 8'h00; 14'h331A: rddata <= 8'h1C; 14'h331B: rddata <= 8'h20;
            14'h331C: rddata <= 8'h20; 14'h331D: rddata <= 8'h20; 14'h331E: rddata <= 8'h1C; 14'h331F: rddata <= 8'h00;
            14'h3320: rddata <= 8'h04; 14'h3321: rddata <= 8'h04; 14'h3322: rddata <= 8'h34; 14'h3323: rddata <= 8'h4C;
            14'h3324: rddata <= 8'h44; 14'h3325: rddata <= 8'h4C; 14'h3326: rddata <= 8'h34; 14'h3327: rddata <= 8'h00;
            14'h3328: rddata <= 8'h00; 14'h3329: rddata <= 8'h00; 14'h332A: rddata <= 8'h38; 14'h332B: rddata <= 8'h44;
            14'h332C: rddata <= 8'h7C; 14'h332D: rddata <= 8'h40; 14'h332E: rddata <= 8'h38; 14'h332F: rddata <= 8'h00;
            14'h3330: rddata <= 8'h08; 14'h3331: rddata <= 8'h10; 14'h3332: rddata <= 8'h10; 14'h3333: rddata <= 8'h38;
            14'h3334: rddata <= 8'h10; 14'h3335: rddata <= 8'h10; 14'h3336: rddata <= 8'h10; 14'h3337: rddata <= 8'h00;
            14'h3338: rddata <= 8'h00; 14'h3339: rddata <= 8'h00; 14'h333A: rddata <= 8'h34; 14'h333B: rddata <= 8'h4C;
            14'h333C: rddata <= 8'h44; 14'h333D: rddata <= 8'h3C; 14'h333E: rddata <= 8'h04; 14'h333F: rddata <= 8'h38;
            14'h3340: rddata <= 8'h40; 14'h3341: rddata <= 8'h40; 14'h3342: rddata <= 8'h78; 14'h3343: rddata <= 8'h44;
            14'h3344: rddata <= 8'h44; 14'h3345: rddata <= 8'h44; 14'h3346: rddata <= 8'h44; 14'h3347: rddata <= 8'h00;
            14'h3348: rddata <= 8'h10; 14'h3349: rddata <= 8'h00; 14'h334A: rddata <= 8'h30; 14'h334B: rddata <= 8'h10;
            14'h334C: rddata <= 8'h10; 14'h334D: rddata <= 8'h10; 14'h334E: rddata <= 8'h38; 14'h334F: rddata <= 8'h00;
            14'h3350: rddata <= 8'h08; 14'h3351: rddata <= 8'h00; 14'h3352: rddata <= 8'h08; 14'h3353: rddata <= 8'h08;
            14'h3354: rddata <= 8'h08; 14'h3355: rddata <= 8'h08; 14'h3356: rddata <= 8'h08; 14'h3357: rddata <= 8'h30;
            14'h3358: rddata <= 8'h40; 14'h3359: rddata <= 8'h40; 14'h335A: rddata <= 8'h48; 14'h335B: rddata <= 8'h50;
            14'h335C: rddata <= 8'h70; 14'h335D: rddata <= 8'h48; 14'h335E: rddata <= 8'h44; 14'h335F: rddata <= 8'h00;
            14'h3360: rddata <= 8'h30; 14'h3361: rddata <= 8'h10; 14'h3362: rddata <= 8'h10; 14'h3363: rddata <= 8'h10;
            14'h3364: rddata <= 8'h10; 14'h3365: rddata <= 8'h10; 14'h3366: rddata <= 8'h38; 14'h3367: rddata <= 8'h00;
            14'h3368: rddata <= 8'h00; 14'h3369: rddata <= 8'h00; 14'h336A: rddata <= 8'h6C; 14'h336B: rddata <= 8'h52;
            14'h336C: rddata <= 8'h52; 14'h336D: rddata <= 8'h52; 14'h336E: rddata <= 8'h52; 14'h336F: rddata <= 8'h00;
            14'h3370: rddata <= 8'h00; 14'h3371: rddata <= 8'h00; 14'h3372: rddata <= 8'h78; 14'h3373: rddata <= 8'h44;
            14'h3374: rddata <= 8'h44; 14'h3375: rddata <= 8'h44; 14'h3376: rddata <= 8'h44; 14'h3377: rddata <= 8'h00;
            14'h3378: rddata <= 8'h00; 14'h3379: rddata <= 8'h00; 14'h337A: rddata <= 8'h38; 14'h337B: rddata <= 8'h44;
            14'h337C: rddata <= 8'h44; 14'h337D: rddata <= 8'h44; 14'h337E: rddata <= 8'h38; 14'h337F: rddata <= 8'h00;
            14'h3380: rddata <= 8'h00; 14'h3381: rddata <= 8'h00; 14'h3382: rddata <= 8'h58; 14'h3383: rddata <= 8'h64;
            14'h3384: rddata <= 8'h44; 14'h3385: rddata <= 8'h64; 14'h3386: rddata <= 8'h58; 14'h3387: rddata <= 8'h40;
            14'h3388: rddata <= 8'h00; 14'h3389: rddata <= 8'h00; 14'h338A: rddata <= 8'h34; 14'h338B: rddata <= 8'h4C;
            14'h338C: rddata <= 8'h44; 14'h338D: rddata <= 8'h4C; 14'h338E: rddata <= 8'h34; 14'h338F: rddata <= 8'h06;
            14'h3390: rddata <= 8'h00; 14'h3391: rddata <= 8'h00; 14'h3392: rddata <= 8'h58; 14'h3393: rddata <= 8'h60;
            14'h3394: rddata <= 8'h40; 14'h3395: rddata <= 8'h40; 14'h3396: rddata <= 8'h40; 14'h3397: rddata <= 8'h00;
            14'h3398: rddata <= 8'h00; 14'h3399: rddata <= 8'h00; 14'h339A: rddata <= 8'h3C; 14'h339B: rddata <= 8'h40;
            14'h339C: rddata <= 8'h38; 14'h339D: rddata <= 8'h04; 14'h339E: rddata <= 8'h78; 14'h339F: rddata <= 8'h00;
            14'h33A0: rddata <= 8'h10; 14'h33A1: rddata <= 8'h10; 14'h33A2: rddata <= 8'h7C; 14'h33A3: rddata <= 8'h10;
            14'h33A4: rddata <= 8'h10; 14'h33A5: rddata <= 8'h10; 14'h33A6: rddata <= 8'h10; 14'h33A7: rddata <= 8'h00;
            14'h33A8: rddata <= 8'h00; 14'h33A9: rddata <= 8'h00; 14'h33AA: rddata <= 8'h44; 14'h33AB: rddata <= 8'h44;
            14'h33AC: rddata <= 8'h44; 14'h33AD: rddata <= 8'h44; 14'h33AE: rddata <= 8'h3C; 14'h33AF: rddata <= 8'h00;
            14'h33B0: rddata <= 8'h00; 14'h33B1: rddata <= 8'h00; 14'h33B2: rddata <= 8'h44; 14'h33B3: rddata <= 8'h44;
            14'h33B4: rddata <= 8'h28; 14'h33B5: rddata <= 8'h28; 14'h33B6: rddata <= 8'h10; 14'h33B7: rddata <= 8'h00;
            14'h33B8: rddata <= 8'h00; 14'h33B9: rddata <= 8'h00; 14'h33BA: rddata <= 8'h52; 14'h33BB: rddata <= 8'h52;
            14'h33BC: rddata <= 8'h52; 14'h33BD: rddata <= 8'h52; 14'h33BE: rddata <= 8'h2C; 14'h33BF: rddata <= 8'h00;
            14'h33C0: rddata <= 8'h00; 14'h33C1: rddata <= 8'h00; 14'h33C2: rddata <= 8'h44; 14'h33C3: rddata <= 8'h28;
            14'h33C4: rddata <= 8'h10; 14'h33C5: rddata <= 8'h28; 14'h33C6: rddata <= 8'h44; 14'h33C7: rddata <= 8'h00;
            14'h33C8: rddata <= 8'h00; 14'h33C9: rddata <= 8'h00; 14'h33CA: rddata <= 8'h24; 14'h33CB: rddata <= 8'h24;
            14'h33CC: rddata <= 8'h24; 14'h33CD: rddata <= 8'h3C; 14'h33CE: rddata <= 8'h04; 14'h33CF: rddata <= 8'h38;
            14'h33D0: rddata <= 8'h00; 14'h33D1: rddata <= 8'h00; 14'h33D2: rddata <= 8'h7C; 14'h33D3: rddata <= 8'h08;
            14'h33D4: rddata <= 8'h10; 14'h33D5: rddata <= 8'h20; 14'h33D6: rddata <= 8'h7C; 14'h33D7: rddata <= 8'h00;
            14'h33D8: rddata <= 8'h0C; 14'h33D9: rddata <= 8'h10; 14'h33DA: rddata <= 8'h10; 14'h33DB: rddata <= 8'h20;
            14'h33DC: rddata <= 8'h10; 14'h33DD: rddata <= 8'h10; 14'h33DE: rddata <= 8'h0C; 14'h33DF: rddata <= 8'h00;
            14'h33E0: rddata <= 8'h10; 14'h33E1: rddata <= 8'h10; 14'h33E2: rddata <= 8'h10; 14'h33E3: rddata <= 8'h00;
            14'h33E4: rddata <= 8'h10; 14'h33E5: rddata <= 8'h10; 14'h33E6: rddata <= 8'h10; 14'h33E7: rddata <= 8'h00;
            14'h33E8: rddata <= 8'h60; 14'h33E9: rddata <= 8'h10; 14'h33EA: rddata <= 8'h10; 14'h33EB: rddata <= 8'h08;
            14'h33EC: rddata <= 8'h10; 14'h33ED: rddata <= 8'h10; 14'h33EE: rddata <= 8'h60; 14'h33EF: rddata <= 8'h00;
            14'h33F0: rddata <= 8'h00; 14'h33F1: rddata <= 8'h00; 14'h33F2: rddata <= 8'h04; 14'h33F3: rddata <= 8'h38;
            14'h33F4: rddata <= 8'h40; 14'h33F5: rddata <= 8'h00; 14'h33F6: rddata <= 8'h00; 14'h33F7: rddata <= 8'h00;
            14'h33F8: rddata <= 8'hFF; 14'h33F9: rddata <= 8'hFF; 14'h33FA: rddata <= 8'hFF; 14'h33FB: rddata <= 8'hFF;
            14'h33FC: rddata <= 8'hFF; 14'h33FD: rddata <= 8'hFF; 14'h33FE: rddata <= 8'hFF; 14'h33FF: rddata <= 8'hFF;
            14'h3400: rddata <= 8'h00; 14'h3401: rddata <= 8'hFF; 14'h3402: rddata <= 8'hFF; 14'h3403: rddata <= 8'hFF;
            14'h3404: rddata <= 8'hFF; 14'h3405: rddata <= 8'hFF; 14'h3406: rddata <= 8'hFF; 14'h3407: rddata <= 8'hFF;
            14'h3408: rddata <= 8'h80; 14'h3409: rddata <= 8'h80; 14'h340A: rddata <= 8'h80; 14'h340B: rddata <= 8'h80;
            14'h340C: rddata <= 8'h80; 14'h340D: rddata <= 8'h80; 14'h340E: rddata <= 8'h80; 14'h340F: rddata <= 8'h80;
            14'h3410: rddata <= 8'h00; 14'h3411: rddata <= 8'h1C; 14'h3412: rddata <= 8'h3C; 14'h3413: rddata <= 8'h00;
            14'h3414: rddata <= 8'h1C; 14'h3415: rddata <= 8'h1E; 14'h3416: rddata <= 8'h3E; 14'h3417: rddata <= 8'hFE;
            14'h3418: rddata <= 8'h3E; 14'h3419: rddata <= 8'h7C; 14'h341A: rddata <= 8'hD8; 14'h341B: rddata <= 8'h78;
            14'h341C: rddata <= 8'h38; 14'h341D: rddata <= 8'h18; 14'h341E: rddata <= 8'h1C; 14'h341F: rddata <= 8'h1C;
            14'h3420: rddata <= 8'h00; 14'h3421: rddata <= 8'h00; 14'h3422: rddata <= 8'h00; 14'h3423: rddata <= 8'h00;
            14'h3424: rddata <= 8'hAA; 14'h3425: rddata <= 8'h55; 14'h3426: rddata <= 8'hAA; 14'h3427: rddata <= 8'h55;
            14'h3428: rddata <= 8'hA0; 14'h3429: rddata <= 8'h50; 14'h342A: rddata <= 8'hA0; 14'h342B: rddata <= 8'h50;
            14'h342C: rddata <= 8'hA0; 14'h342D: rddata <= 8'h50; 14'h342E: rddata <= 8'hA0; 14'h342F: rddata <= 8'h50;
            14'h3430: rddata <= 8'hAA; 14'h3431: rddata <= 8'h55; 14'h3432: rddata <= 8'hAA; 14'h3433: rddata <= 8'h55;
            14'h3434: rddata <= 8'hAA; 14'h3435: rddata <= 8'h55; 14'h3436: rddata <= 8'hAA; 14'h3437: rddata <= 8'h55;
            14'h3438: rddata <= 8'h00; 14'h3439: rddata <= 8'h18; 14'h343A: rddata <= 8'h3C; 14'h343B: rddata <= 8'h7E;
            14'h343C: rddata <= 8'h7E; 14'h343D: rddata <= 8'h3C; 14'h343E: rddata <= 8'h18; 14'h343F: rddata <= 8'h00;
            14'h3440: rddata <= 8'h00; 14'h3441: rddata <= 8'h00; 14'h3442: rddata <= 8'h00; 14'h3443: rddata <= 8'h00;
            14'h3444: rddata <= 8'h00; 14'h3445: rddata <= 8'h00; 14'h3446: rddata <= 8'hFF; 14'h3447: rddata <= 8'hFF;
            14'h3448: rddata <= 8'h00; 14'h3449: rddata <= 8'h00; 14'h344A: rddata <= 8'hFF; 14'h344B: rddata <= 8'hFF;
            14'h344C: rddata <= 8'hFF; 14'h344D: rddata <= 8'hFF; 14'h344E: rddata <= 8'hFF; 14'h344F: rddata <= 8'hFF;
            14'h3450: rddata <= 8'h18; 14'h3451: rddata <= 8'h18; 14'h3452: rddata <= 8'h3C; 14'h3453: rddata <= 8'h7E;
            14'h3454: rddata <= 8'hFF; 14'h3455: rddata <= 8'hDB; 14'h3456: rddata <= 8'h18; 14'h3457: rddata <= 8'h3C;
            14'h3458: rddata <= 8'h3C; 14'h3459: rddata <= 8'h18; 14'h345A: rddata <= 8'hDB; 14'h345B: rddata <= 8'hFF;
            14'h345C: rddata <= 8'h7E; 14'h345D: rddata <= 8'h3C; 14'h345E: rddata <= 8'h18; 14'h345F: rddata <= 8'h18;
            14'h3460: rddata <= 8'h00; 14'h3461: rddata <= 8'h1C; 14'h3462: rddata <= 8'h3C; 14'h3463: rddata <= 8'h00;
            14'h3464: rddata <= 8'h9C; 14'h3465: rddata <= 8'h9E; 14'h3466: rddata <= 8'hFB; 14'h3467: rddata <= 8'h3B;
            14'h3468: rddata <= 8'h3E; 14'h3469: rddata <= 8'hFC; 14'h346A: rddata <= 8'hF8; 14'h346B: rddata <= 8'hDC;
            14'h346C: rddata <= 8'hCF; 14'h346D: rddata <= 8'hC3; 14'h346E: rddata <= 8'h01; 14'h346F: rddata <= 8'h00;
            14'h3470: rddata <= 8'hC0; 14'h3471: rddata <= 8'hF0; 14'h3472: rddata <= 8'hFC; 14'h3473: rddata <= 8'hFF;
            14'h3474: rddata <= 8'hFF; 14'h3475: rddata <= 8'hFC; 14'h3476: rddata <= 8'hF0; 14'h3477: rddata <= 8'hC0;
            14'h3478: rddata <= 8'h18; 14'h3479: rddata <= 8'h18; 14'h347A: rddata <= 8'h3C; 14'h347B: rddata <= 8'h3C;
            14'h347C: rddata <= 8'h7E; 14'h347D: rddata <= 8'h7E; 14'h347E: rddata <= 8'hFF; 14'h347F: rddata <= 8'hFF;
            14'h3480: rddata <= 8'h00; 14'h3481: rddata <= 8'h00; 14'h3482: rddata <= 8'h00; 14'h3483: rddata <= 8'h00;
            14'h3484: rddata <= 8'h00; 14'h3485: rddata <= 8'h00; 14'h3486: rddata <= 8'h00; 14'h3487: rddata <= 8'hFF;
            14'h3488: rddata <= 8'hFE; 14'h3489: rddata <= 8'hFE; 14'h348A: rddata <= 8'hFE; 14'h348B: rddata <= 8'hFE;
            14'h348C: rddata <= 8'hFE; 14'h348D: rddata <= 8'hFE; 14'h348E: rddata <= 8'hFE; 14'h348F: rddata <= 8'hFE;
            14'h3490: rddata <= 8'h3C; 14'h3491: rddata <= 8'h52; 14'h3492: rddata <= 8'h3C; 14'h3493: rddata <= 8'h80;
            14'h3494: rddata <= 8'hBC; 14'h3495: rddata <= 8'hFF; 14'h3496: rddata <= 8'h3D; 14'h3497: rddata <= 8'h3D;
            14'h3498: rddata <= 8'h3C; 14'h3499: rddata <= 8'h4A; 14'h349A: rddata <= 8'h3C; 14'h349B: rddata <= 8'h01;
            14'h349C: rddata <= 8'h3D; 14'h349D: rddata <= 8'hFF; 14'h349E: rddata <= 8'hBC; 14'h349F: rddata <= 8'hBC;
            14'h34A0: rddata <= 8'hAA; 14'h34A1: rddata <= 8'h55; 14'h34A2: rddata <= 8'hAA; 14'h34A3: rddata <= 8'h55;
            14'h34A4: rddata <= 8'h00; 14'h34A5: rddata <= 8'h00; 14'h34A6: rddata <= 8'h00; 14'h34A7: rddata <= 8'h00;
            14'h34A8: rddata <= 8'h0A; 14'h34A9: rddata <= 8'h05; 14'h34AA: rddata <= 8'h0A; 14'h34AB: rddata <= 8'h05;
            14'h34AC: rddata <= 8'h0A; 14'h34AD: rddata <= 8'h05; 14'h34AE: rddata <= 8'h0A; 14'h34AF: rddata <= 8'h05;
            14'h34B0: rddata <= 8'h3C; 14'h34B1: rddata <= 8'h7E; 14'h34B2: rddata <= 8'hFF; 14'h34B3: rddata <= 8'hFF;
            14'h34B4: rddata <= 8'hFF; 14'h34B5: rddata <= 8'hFF; 14'h34B6: rddata <= 8'h7E; 14'h34B7: rddata <= 8'h3C;
            14'h34B8: rddata <= 8'hC0; 14'h34B9: rddata <= 8'hC0; 14'h34BA: rddata <= 8'hC0; 14'h34BB: rddata <= 8'hC0;
            14'h34BC: rddata <= 8'hC0; 14'h34BD: rddata <= 8'hC0; 14'h34BE: rddata <= 8'hC0; 14'h34BF: rddata <= 8'hC0;
            14'h34C0: rddata <= 8'hE0; 14'h34C1: rddata <= 8'hE0; 14'h34C2: rddata <= 8'hE0; 14'h34C3: rddata <= 8'hE0;
            14'h34C4: rddata <= 8'hE0; 14'h34C5: rddata <= 8'hE0; 14'h34C6: rddata <= 8'hE0; 14'h34C7: rddata <= 8'hE0;
            14'h34C8: rddata <= 8'hF8; 14'h34C9: rddata <= 8'hF8; 14'h34CA: rddata <= 8'hF8; 14'h34CB: rddata <= 8'hF8;
            14'h34CC: rddata <= 8'hF8; 14'h34CD: rddata <= 8'hF8; 14'h34CE: rddata <= 8'hF8; 14'h34CF: rddata <= 8'hF8;
            14'h34D0: rddata <= 8'h30; 14'h34D1: rddata <= 8'h38; 14'h34D2: rddata <= 8'h9C; 14'h34D3: rddata <= 8'hFF;
            14'h34D4: rddata <= 8'hFF; 14'h34D5: rddata <= 8'h9C; 14'h34D6: rddata <= 8'h38; 14'h34D7: rddata <= 8'h30;
            14'h34D8: rddata <= 8'h0C; 14'h34D9: rddata <= 8'h1C; 14'h34DA: rddata <= 8'h39; 14'h34DB: rddata <= 8'hFF;
            14'h34DC: rddata <= 8'hFF; 14'h34DD: rddata <= 8'h39; 14'h34DE: rddata <= 8'h1C; 14'h34DF: rddata <= 8'h0C;
            14'h34E0: rddata <= 8'h00; 14'h34E1: rddata <= 8'h66; 14'h34E2: rddata <= 8'h7E; 14'h34E3: rddata <= 8'h42;
            14'h34E4: rddata <= 8'hC3; 14'h34E5: rddata <= 8'hFF; 14'h34E6: rddata <= 8'h18; 14'h34E7: rddata <= 8'h00;
            14'h34E8: rddata <= 8'h00; 14'h34E9: rddata <= 8'h18; 14'h34EA: rddata <= 8'hFF; 14'h34EB: rddata <= 8'hC3;
            14'h34EC: rddata <= 8'h42; 14'h34ED: rddata <= 8'h7E; 14'h34EE: rddata <= 8'h66; 14'h34EF: rddata <= 8'h00;
            14'h34F0: rddata <= 8'h03; 14'h34F1: rddata <= 8'h0F; 14'h34F2: rddata <= 8'h3F; 14'h34F3: rddata <= 8'hFF;
            14'h34F4: rddata <= 8'hFF; 14'h34F5: rddata <= 8'h3F; 14'h34F6: rddata <= 8'h0F; 14'h34F7: rddata <= 8'h03;
            14'h34F8: rddata <= 8'hFF; 14'h34F9: rddata <= 8'hFF; 14'h34FA: rddata <= 8'h7E; 14'h34FB: rddata <= 8'h7E;
            14'h34FC: rddata <= 8'h3C; 14'h34FD: rddata <= 8'h3C; 14'h34FE: rddata <= 8'h18; 14'h34FF: rddata <= 8'h18;
            14'h3500: rddata <= 8'h00; 14'h3501: rddata <= 8'h00; 14'h3502: rddata <= 8'h00; 14'h3503: rddata <= 8'h00;
            14'h3504: rddata <= 8'h00; 14'h3505: rddata <= 8'h00; 14'h3506: rddata <= 8'h00; 14'h3507: rddata <= 8'h00;
            14'h3508: rddata <= 8'hF0; 14'h3509: rddata <= 8'hF0; 14'h350A: rddata <= 8'hF0; 14'h350B: rddata <= 8'h00;
            14'h350C: rddata <= 8'h00; 14'h350D: rddata <= 8'h00; 14'h350E: rddata <= 8'h00; 14'h350F: rddata <= 8'h00;
            14'h3510: rddata <= 8'h0F; 14'h3511: rddata <= 8'h0F; 14'h3512: rddata <= 8'h0F; 14'h3513: rddata <= 8'h00;
            14'h3514: rddata <= 8'h00; 14'h3515: rddata <= 8'h00; 14'h3516: rddata <= 8'h00; 14'h3517: rddata <= 8'h00;
            14'h3518: rddata <= 8'hFF; 14'h3519: rddata <= 8'hFF; 14'h351A: rddata <= 8'hFF; 14'h351B: rddata <= 8'h00;
            14'h351C: rddata <= 8'h00; 14'h351D: rddata <= 8'h00; 14'h351E: rddata <= 8'h00; 14'h351F: rddata <= 8'h00;
            14'h3520: rddata <= 8'h00; 14'h3521: rddata <= 8'h00; 14'h3522: rddata <= 8'h00; 14'h3523: rddata <= 8'hF0;
            14'h3524: rddata <= 8'hF0; 14'h3525: rddata <= 8'h00; 14'h3526: rddata <= 8'h00; 14'h3527: rddata <= 8'h00;
            14'h3528: rddata <= 8'hF0; 14'h3529: rddata <= 8'hF0; 14'h352A: rddata <= 8'hF0; 14'h352B: rddata <= 8'hF0;
            14'h352C: rddata <= 8'hF0; 14'h352D: rddata <= 8'h00; 14'h352E: rddata <= 8'h00; 14'h352F: rddata <= 8'h00;
            14'h3530: rddata <= 8'h0F; 14'h3531: rddata <= 8'h0F; 14'h3532: rddata <= 8'h0F; 14'h3533: rddata <= 8'hF0;
            14'h3534: rddata <= 8'hF0; 14'h3535: rddata <= 8'h00; 14'h3536: rddata <= 8'h00; 14'h3537: rddata <= 8'h00;
            14'h3538: rddata <= 8'hFF; 14'h3539: rddata <= 8'hFF; 14'h353A: rddata <= 8'hFF; 14'h353B: rddata <= 8'hF0;
            14'h353C: rddata <= 8'hF0; 14'h353D: rddata <= 8'h00; 14'h353E: rddata <= 8'h00; 14'h353F: rddata <= 8'h00;
            14'h3540: rddata <= 8'h00; 14'h3541: rddata <= 8'h00; 14'h3542: rddata <= 8'h00; 14'h3543: rddata <= 8'h0F;
            14'h3544: rddata <= 8'h0F; 14'h3545: rddata <= 8'h00; 14'h3546: rddata <= 8'h00; 14'h3547: rddata <= 8'h00;
            14'h3548: rddata <= 8'hF0; 14'h3549: rddata <= 8'hF0; 14'h354A: rddata <= 8'hF0; 14'h354B: rddata <= 8'h0F;
            14'h354C: rddata <= 8'h0F; 14'h354D: rddata <= 8'h00; 14'h354E: rddata <= 8'h00; 14'h354F: rddata <= 8'h00;
            14'h3550: rddata <= 8'h0F; 14'h3551: rddata <= 8'h0F; 14'h3552: rddata <= 8'h0F; 14'h3553: rddata <= 8'h0F;
            14'h3554: rddata <= 8'h0F; 14'h3555: rddata <= 8'h00; 14'h3556: rddata <= 8'h00; 14'h3557: rddata <= 8'h00;
            14'h3558: rddata <= 8'hFF; 14'h3559: rddata <= 8'hFF; 14'h355A: rddata <= 8'hFF; 14'h355B: rddata <= 8'h0F;
            14'h355C: rddata <= 8'h0F; 14'h355D: rddata <= 8'h00; 14'h355E: rddata <= 8'h00; 14'h355F: rddata <= 8'h00;
            14'h3560: rddata <= 8'h00; 14'h3561: rddata <= 8'h00; 14'h3562: rddata <= 8'h00; 14'h3563: rddata <= 8'hFF;
            14'h3564: rddata <= 8'hFF; 14'h3565: rddata <= 8'h00; 14'h3566: rddata <= 8'h00; 14'h3567: rddata <= 8'h00;
            14'h3568: rddata <= 8'hF0; 14'h3569: rddata <= 8'hF0; 14'h356A: rddata <= 8'hF0; 14'h356B: rddata <= 8'hFF;
            14'h356C: rddata <= 8'hFF; 14'h356D: rddata <= 8'h00; 14'h356E: rddata <= 8'h00; 14'h356F: rddata <= 8'h00;
            14'h3570: rddata <= 8'h0F; 14'h3571: rddata <= 8'h0F; 14'h3572: rddata <= 8'h0F; 14'h3573: rddata <= 8'hFF;
            14'h3574: rddata <= 8'hFF; 14'h3575: rddata <= 8'h00; 14'h3576: rddata <= 8'h00; 14'h3577: rddata <= 8'h00;
            14'h3578: rddata <= 8'hFF; 14'h3579: rddata <= 8'hFF; 14'h357A: rddata <= 8'hFF; 14'h357B: rddata <= 8'hFF;
            14'h357C: rddata <= 8'hFF; 14'h357D: rddata <= 8'h00; 14'h357E: rddata <= 8'h00; 14'h357F: rddata <= 8'h00;
            14'h3580: rddata <= 8'h00; 14'h3581: rddata <= 8'h00; 14'h3582: rddata <= 8'h00; 14'h3583: rddata <= 8'h00;
            14'h3584: rddata <= 8'h00; 14'h3585: rddata <= 8'hF0; 14'h3586: rddata <= 8'hF0; 14'h3587: rddata <= 8'hF0;
            14'h3588: rddata <= 8'hF0; 14'h3589: rddata <= 8'hF0; 14'h358A: rddata <= 8'hF0; 14'h358B: rddata <= 8'h00;
            14'h358C: rddata <= 8'h00; 14'h358D: rddata <= 8'hF0; 14'h358E: rddata <= 8'hF0; 14'h358F: rddata <= 8'hF0;
            14'h3590: rddata <= 8'h0F; 14'h3591: rddata <= 8'h0F; 14'h3592: rddata <= 8'h0F; 14'h3593: rddata <= 8'h00;
            14'h3594: rddata <= 8'h00; 14'h3595: rddata <= 8'hF0; 14'h3596: rddata <= 8'hF0; 14'h3597: rddata <= 8'hF0;
            14'h3598: rddata <= 8'hFF; 14'h3599: rddata <= 8'hFF; 14'h359A: rddata <= 8'hFF; 14'h359B: rddata <= 8'h00;
            14'h359C: rddata <= 8'h00; 14'h359D: rddata <= 8'hF0; 14'h359E: rddata <= 8'hF0; 14'h359F: rddata <= 8'hF0;
            14'h35A0: rddata <= 8'h00; 14'h35A1: rddata <= 8'h00; 14'h35A2: rddata <= 8'h00; 14'h35A3: rddata <= 8'hF0;
            14'h35A4: rddata <= 8'hF0; 14'h35A5: rddata <= 8'hF0; 14'h35A6: rddata <= 8'hF0; 14'h35A7: rddata <= 8'hF0;
            14'h35A8: rddata <= 8'hF0; 14'h35A9: rddata <= 8'hF0; 14'h35AA: rddata <= 8'hF0; 14'h35AB: rddata <= 8'hF0;
            14'h35AC: rddata <= 8'hF0; 14'h35AD: rddata <= 8'hF0; 14'h35AE: rddata <= 8'hF0; 14'h35AF: rddata <= 8'hF0;
            14'h35B0: rddata <= 8'h0F; 14'h35B1: rddata <= 8'h0F; 14'h35B2: rddata <= 8'h0F; 14'h35B3: rddata <= 8'hF0;
            14'h35B4: rddata <= 8'hF0; 14'h35B5: rddata <= 8'hF0; 14'h35B6: rddata <= 8'hF0; 14'h35B7: rddata <= 8'hF0;
            14'h35B8: rddata <= 8'hFF; 14'h35B9: rddata <= 8'hFF; 14'h35BA: rddata <= 8'hFF; 14'h35BB: rddata <= 8'hF0;
            14'h35BC: rddata <= 8'hF0; 14'h35BD: rddata <= 8'hF0; 14'h35BE: rddata <= 8'hF0; 14'h35BF: rddata <= 8'hF0;
            14'h35C0: rddata <= 8'h00; 14'h35C1: rddata <= 8'h00; 14'h35C2: rddata <= 8'h00; 14'h35C3: rddata <= 8'h0F;
            14'h35C4: rddata <= 8'h0F; 14'h35C5: rddata <= 8'hF0; 14'h35C6: rddata <= 8'hF0; 14'h35C7: rddata <= 8'hF0;
            14'h35C8: rddata <= 8'hF0; 14'h35C9: rddata <= 8'hF0; 14'h35CA: rddata <= 8'hF0; 14'h35CB: rddata <= 8'h0F;
            14'h35CC: rddata <= 8'h0F; 14'h35CD: rddata <= 8'hF0; 14'h35CE: rddata <= 8'hF0; 14'h35CF: rddata <= 8'hF0;
            14'h35D0: rddata <= 8'h0F; 14'h35D1: rddata <= 8'h0F; 14'h35D2: rddata <= 8'h0F; 14'h35D3: rddata <= 8'h0F;
            14'h35D4: rddata <= 8'h0F; 14'h35D5: rddata <= 8'hF0; 14'h35D6: rddata <= 8'hF0; 14'h35D7: rddata <= 8'hF0;
            14'h35D8: rddata <= 8'hFF; 14'h35D9: rddata <= 8'hFF; 14'h35DA: rddata <= 8'hFF; 14'h35DB: rddata <= 8'h0F;
            14'h35DC: rddata <= 8'h0F; 14'h35DD: rddata <= 8'hF0; 14'h35DE: rddata <= 8'hF0; 14'h35DF: rddata <= 8'hF0;
            14'h35E0: rddata <= 8'h00; 14'h35E1: rddata <= 8'h00; 14'h35E2: rddata <= 8'h00; 14'h35E3: rddata <= 8'hFF;
            14'h35E4: rddata <= 8'hFF; 14'h35E5: rddata <= 8'hF0; 14'h35E6: rddata <= 8'hF0; 14'h35E7: rddata <= 8'hF0;
            14'h35E8: rddata <= 8'hF0; 14'h35E9: rddata <= 8'hF0; 14'h35EA: rddata <= 8'hF0; 14'h35EB: rddata <= 8'hFF;
            14'h35EC: rddata <= 8'hFF; 14'h35ED: rddata <= 8'hF0; 14'h35EE: rddata <= 8'hF0; 14'h35EF: rddata <= 8'hF0;
            14'h35F0: rddata <= 8'h0F; 14'h35F1: rddata <= 8'h0F; 14'h35F2: rddata <= 8'h0F; 14'h35F3: rddata <= 8'hFF;
            14'h35F4: rddata <= 8'hFF; 14'h35F5: rddata <= 8'hF0; 14'h35F6: rddata <= 8'hF0; 14'h35F7: rddata <= 8'hF0;
            14'h35F8: rddata <= 8'hFF; 14'h35F9: rddata <= 8'hFF; 14'h35FA: rddata <= 8'hFF; 14'h35FB: rddata <= 8'hFF;
            14'h35FC: rddata <= 8'hFF; 14'h35FD: rddata <= 8'hF0; 14'h35FE: rddata <= 8'hF0; 14'h35FF: rddata <= 8'hF0;
            14'h3600: rddata <= 8'h01; 14'h3601: rddata <= 8'h03; 14'h3602: rddata <= 8'h07; 14'h3603: rddata <= 8'h0F;
            14'h3604: rddata <= 8'h1F; 14'h3605: rddata <= 8'h3F; 14'h3606: rddata <= 8'h7F; 14'h3607: rddata <= 8'hFF;
            14'h3608: rddata <= 8'h80; 14'h3609: rddata <= 8'hC0; 14'h360A: rddata <= 8'hE0; 14'h360B: rddata <= 8'hF0;
            14'h360C: rddata <= 8'hF8; 14'h360D: rddata <= 8'hFC; 14'h360E: rddata <= 8'hFE; 14'h360F: rddata <= 8'hFF;
            14'h3610: rddata <= 8'hFF; 14'h3611: rddata <= 8'hFF; 14'h3612: rddata <= 8'h7E; 14'h3613: rddata <= 8'h3C;
            14'h3614: rddata <= 8'h00; 14'h3615: rddata <= 8'h00; 14'h3616: rddata <= 8'h00; 14'h3617: rddata <= 8'h00;
            14'h3618: rddata <= 8'hFC; 14'h3619: rddata <= 8'hFC; 14'h361A: rddata <= 8'hFC; 14'h361B: rddata <= 8'hFC;
            14'h361C: rddata <= 8'hFC; 14'h361D: rddata <= 8'hFC; 14'h361E: rddata <= 8'hFC; 14'h361F: rddata <= 8'hFC;
            14'h3620: rddata <= 8'h00; 14'h3621: rddata <= 8'h00; 14'h3622: rddata <= 8'h3C; 14'h3623: rddata <= 8'h3C;
            14'h3624: rddata <= 8'h3C; 14'h3625: rddata <= 8'h3C; 14'h3626: rddata <= 8'h00; 14'h3627: rddata <= 8'h00;
            14'h3628: rddata <= 8'h18; 14'h3629: rddata <= 8'h3C; 14'h362A: rddata <= 8'h7E; 14'h362B: rddata <= 8'hFF;
            14'h362C: rddata <= 8'hFF; 14'h362D: rddata <= 8'h7E; 14'h362E: rddata <= 8'h3C; 14'h362F: rddata <= 8'h18;
            14'h3630: rddata <= 8'h00; 14'h3631: rddata <= 8'h00; 14'h3632: rddata <= 8'h00; 14'h3633: rddata <= 8'h18;
            14'h3634: rddata <= 8'h18; 14'h3635: rddata <= 8'h00; 14'h3636: rddata <= 8'h00; 14'h3637: rddata <= 8'h00;
            14'h3638: rddata <= 8'h0F; 14'h3639: rddata <= 8'h0F; 14'h363A: rddata <= 8'h07; 14'h363B: rddata <= 8'h03;
            14'h363C: rddata <= 8'h00; 14'h363D: rddata <= 8'h00; 14'h363E: rddata <= 8'h00; 14'h363F: rddata <= 8'h00;
            14'h3640: rddata <= 8'h18; 14'h3641: rddata <= 8'h18; 14'h3642: rddata <= 8'h18; 14'h3643: rddata <= 8'hFF;
            14'h3644: rddata <= 8'hFF; 14'h3645: rddata <= 8'h18; 14'h3646: rddata <= 8'h18; 14'h3647: rddata <= 8'h18;
            14'h3648: rddata <= 8'h00; 14'h3649: rddata <= 8'h00; 14'h364A: rddata <= 8'h00; 14'h364B: rddata <= 8'h00;
            14'h364C: rddata <= 8'hC0; 14'h364D: rddata <= 8'hE0; 14'h364E: rddata <= 8'hF0; 14'h364F: rddata <= 8'hF0;
            14'h3650: rddata <= 8'h01; 14'h3651: rddata <= 8'h02; 14'h3652: rddata <= 8'h04; 14'h3653: rddata <= 8'h08;
            14'h3654: rddata <= 8'h10; 14'h3655: rddata <= 8'h20; 14'h3656: rddata <= 8'h40; 14'h3657: rddata <= 8'h80;
            14'h3658: rddata <= 8'h03; 14'h3659: rddata <= 8'h07; 14'h365A: rddata <= 8'h0F; 14'h365B: rddata <= 8'h0F;
            14'h365C: rddata <= 8'h0F; 14'h365D: rddata <= 8'h0F; 14'h365E: rddata <= 8'h07; 14'h365F: rddata <= 8'h03;
            14'h3660: rddata <= 8'h18; 14'h3661: rddata <= 8'h18; 14'h3662: rddata <= 8'h18; 14'h3663: rddata <= 8'hFF;
            14'h3664: rddata <= 8'hFF; 14'h3665: rddata <= 8'h00; 14'h3666: rddata <= 8'h00; 14'h3667: rddata <= 8'h00;
            14'h3668: rddata <= 8'h18; 14'h3669: rddata <= 8'h18; 14'h366A: rddata <= 8'h18; 14'h366B: rddata <= 8'h1F;
            14'h366C: rddata <= 8'h1F; 14'h366D: rddata <= 8'h18; 14'h366E: rddata <= 8'h18; 14'h366F: rddata <= 8'h18;
            14'h3670: rddata <= 8'h00; 14'h3671: rddata <= 8'h00; 14'h3672: rddata <= 8'h00; 14'h3673: rddata <= 8'hF8;
            14'h3674: rddata <= 8'hF8; 14'h3675: rddata <= 8'h18; 14'h3676: rddata <= 8'h18; 14'h3677: rddata <= 8'h18;
            14'h3678: rddata <= 8'h18; 14'h3679: rddata <= 8'h18; 14'h367A: rddata <= 8'h18; 14'h367B: rddata <= 8'h1F;
            14'h367C: rddata <= 8'h1F; 14'h367D: rddata <= 8'h00; 14'h367E: rddata <= 8'h00; 14'h367F: rddata <= 8'h00;
            14'h3680: rddata <= 8'h09; 14'h3681: rddata <= 8'h20; 14'h3682: rddata <= 8'h04; 14'h3683: rddata <= 8'h80;
            14'h3684: rddata <= 8'h11; 14'h3685: rddata <= 8'h40; 14'h3686: rddata <= 8'h08; 14'h3687: rddata <= 8'h02;
            14'h3688: rddata <= 8'h52; 14'h3689: rddata <= 8'h44; 14'h368A: rddata <= 8'h2D; 14'h368B: rddata <= 8'hC4;
            14'h368C: rddata <= 8'h11; 14'h368D: rddata <= 8'hB4; 14'h368E: rddata <= 8'h23; 14'h368F: rddata <= 8'h4A;
            14'h3690: rddata <= 8'h00; 14'h3691: rddata <= 8'h00; 14'h3692: rddata <= 8'h00; 14'h3693: rddata <= 8'h00;
            14'h3694: rddata <= 8'h3C; 14'h3695: rddata <= 8'h7E; 14'h3696: rddata <= 8'hFF; 14'h3697: rddata <= 8'hFF;
            14'h3698: rddata <= 8'h00; 14'h3699: rddata <= 8'h10; 14'h369A: rddata <= 8'h2C; 14'h369B: rddata <= 8'h3A;
            14'h369C: rddata <= 8'h5C; 14'h369D: rddata <= 8'h34; 14'h369E: rddata <= 8'h04; 14'h369F: rddata <= 8'h00;
            14'h36A0: rddata <= 8'h66; 14'h36A1: rddata <= 8'hFF; 14'h36A2: rddata <= 8'hFF; 14'h36A3: rddata <= 8'hFF;
            14'h36A4: rddata <= 8'h7E; 14'h36A5: rddata <= 8'h3C; 14'h36A6: rddata <= 8'h18; 14'h36A7: rddata <= 8'h18;
            14'h36A8: rddata <= 8'h18; 14'h36A9: rddata <= 8'h3C; 14'h36AA: rddata <= 8'h18; 14'h36AB: rddata <= 8'h42;
            14'h36AC: rddata <= 8'hE7; 14'h36AD: rddata <= 8'h42; 14'h36AE: rddata <= 8'h18; 14'h36AF: rddata <= 8'h3C;
            14'h36B0: rddata <= 8'h18; 14'h36B1: rddata <= 8'h18; 14'h36B2: rddata <= 8'h18; 14'h36B3: rddata <= 8'h18;
            14'h36B4: rddata <= 8'h18; 14'h36B5: rddata <= 8'h18; 14'h36B6: rddata <= 8'h18; 14'h36B7: rddata <= 8'h18;
            14'h36B8: rddata <= 8'h00; 14'h36B9: rddata <= 8'h00; 14'h36BA: rddata <= 8'h00; 14'h36BB: rddata <= 8'h00;
            14'h36BC: rddata <= 8'h03; 14'h36BD: rddata <= 8'h07; 14'h36BE: rddata <= 8'h0F; 14'h36BF: rddata <= 8'h0F;
            14'h36C0: rddata <= 8'h81; 14'h36C1: rddata <= 8'h42; 14'h36C2: rddata <= 8'h24; 14'h36C3: rddata <= 8'h18;
            14'h36C4: rddata <= 8'h18; 14'h36C5: rddata <= 8'h24; 14'h36C6: rddata <= 8'h42; 14'h36C7: rddata <= 8'h81;
            14'h36C8: rddata <= 8'hF0; 14'h36C9: rddata <= 8'hF0; 14'h36CA: rddata <= 8'hE0; 14'h36CB: rddata <= 8'hC0;
            14'h36CC: rddata <= 8'h00; 14'h36CD: rddata <= 8'h00; 14'h36CE: rddata <= 8'h00; 14'h36CF: rddata <= 8'h00;
            14'h36D0: rddata <= 8'h80; 14'h36D1: rddata <= 8'h40; 14'h36D2: rddata <= 8'h20; 14'h36D3: rddata <= 8'h10;
            14'h36D4: rddata <= 8'h08; 14'h36D5: rddata <= 8'h04; 14'h36D6: rddata <= 8'h02; 14'h36D7: rddata <= 8'h01;
            14'h36D8: rddata <= 8'hC0; 14'h36D9: rddata <= 8'hE0; 14'h36DA: rddata <= 8'hF0; 14'h36DB: rddata <= 8'hF0;
            14'h36DC: rddata <= 8'hF0; 14'h36DD: rddata <= 8'hF0; 14'h36DE: rddata <= 8'hE0; 14'h36DF: rddata <= 8'hC0;
            14'h36E0: rddata <= 8'h00; 14'h36E1: rddata <= 8'h00; 14'h36E2: rddata <= 8'h00; 14'h36E3: rddata <= 8'hFF;
            14'h36E4: rddata <= 8'hFF; 14'h36E5: rddata <= 8'h18; 14'h36E6: rddata <= 8'h18; 14'h36E7: rddata <= 8'h18;
            14'h36E8: rddata <= 8'h18; 14'h36E9: rddata <= 8'h18; 14'h36EA: rddata <= 8'h18; 14'h36EB: rddata <= 8'hF8;
            14'h36EC: rddata <= 8'hF8; 14'h36ED: rddata <= 8'h18; 14'h36EE: rddata <= 8'h18; 14'h36EF: rddata <= 8'h18;
            14'h36F0: rddata <= 8'h00; 14'h36F1: rddata <= 8'h00; 14'h36F2: rddata <= 8'h00; 14'h36F3: rddata <= 8'h1F;
            14'h36F4: rddata <= 8'h1F; 14'h36F5: rddata <= 8'h18; 14'h36F6: rddata <= 8'h18; 14'h36F7: rddata <= 8'h18;
            14'h36F8: rddata <= 8'h18; 14'h36F9: rddata <= 8'h18; 14'h36FA: rddata <= 8'h18; 14'h36FB: rddata <= 8'hF8;
            14'h36FC: rddata <= 8'hF8; 14'h36FD: rddata <= 8'h00; 14'h36FE: rddata <= 8'h00; 14'h36FF: rddata <= 8'h00;
            14'h3700: rddata <= 8'h00; 14'h3701: rddata <= 8'h00; 14'h3702: rddata <= 8'h00; 14'h3703: rddata <= 8'h00;
            14'h3704: rddata <= 8'h00; 14'h3705: rddata <= 8'h0F; 14'h3706: rddata <= 8'h0F; 14'h3707: rddata <= 8'h0F;
            14'h3708: rddata <= 8'hF0; 14'h3709: rddata <= 8'hF0; 14'h370A: rddata <= 8'hF0; 14'h370B: rddata <= 8'h00;
            14'h370C: rddata <= 8'h00; 14'h370D: rddata <= 8'h0F; 14'h370E: rddata <= 8'h0F; 14'h370F: rddata <= 8'h0F;
            14'h3710: rddata <= 8'h0F; 14'h3711: rddata <= 8'h0F; 14'h3712: rddata <= 8'h0F; 14'h3713: rddata <= 8'h00;
            14'h3714: rddata <= 8'h00; 14'h3715: rddata <= 8'h0F; 14'h3716: rddata <= 8'h0F; 14'h3717: rddata <= 8'h0F;
            14'h3718: rddata <= 8'hFF; 14'h3719: rddata <= 8'hFF; 14'h371A: rddata <= 8'hFF; 14'h371B: rddata <= 8'h00;
            14'h371C: rddata <= 8'h00; 14'h371D: rddata <= 8'h0F; 14'h371E: rddata <= 8'h0F; 14'h371F: rddata <= 8'h0F;
            14'h3720: rddata <= 8'h00; 14'h3721: rddata <= 8'h00; 14'h3722: rddata <= 8'h00; 14'h3723: rddata <= 8'hF0;
            14'h3724: rddata <= 8'hF0; 14'h3725: rddata <= 8'h0F; 14'h3726: rddata <= 8'h0F; 14'h3727: rddata <= 8'h0F;
            14'h3728: rddata <= 8'hF0; 14'h3729: rddata <= 8'hF0; 14'h372A: rddata <= 8'hF0; 14'h372B: rddata <= 8'hF0;
            14'h372C: rddata <= 8'hF0; 14'h372D: rddata <= 8'h0F; 14'h372E: rddata <= 8'h0F; 14'h372F: rddata <= 8'h0F;
            14'h3730: rddata <= 8'h0F; 14'h3731: rddata <= 8'h0F; 14'h3732: rddata <= 8'h0F; 14'h3733: rddata <= 8'hF0;
            14'h3734: rddata <= 8'hF0; 14'h3735: rddata <= 8'h0F; 14'h3736: rddata <= 8'h0F; 14'h3737: rddata <= 8'h0F;
            14'h3738: rddata <= 8'hFF; 14'h3739: rddata <= 8'hFF; 14'h373A: rddata <= 8'hFF; 14'h373B: rddata <= 8'hF0;
            14'h373C: rddata <= 8'hF0; 14'h373D: rddata <= 8'h0F; 14'h373E: rddata <= 8'h0F; 14'h373F: rddata <= 8'h0F;
            14'h3740: rddata <= 8'h00; 14'h3741: rddata <= 8'h00; 14'h3742: rddata <= 8'h00; 14'h3743: rddata <= 8'h0F;
            14'h3744: rddata <= 8'h0F; 14'h3745: rddata <= 8'h0F; 14'h3746: rddata <= 8'h0F; 14'h3747: rddata <= 8'h0F;
            14'h3748: rddata <= 8'hF0; 14'h3749: rddata <= 8'hF0; 14'h374A: rddata <= 8'hF0; 14'h374B: rddata <= 8'h0F;
            14'h374C: rddata <= 8'h0F; 14'h374D: rddata <= 8'h0F; 14'h374E: rddata <= 8'h0F; 14'h374F: rddata <= 8'h0F;
            14'h3750: rddata <= 8'h0F; 14'h3751: rddata <= 8'h0F; 14'h3752: rddata <= 8'h0F; 14'h3753: rddata <= 8'h0F;
            14'h3754: rddata <= 8'h0F; 14'h3755: rddata <= 8'h0F; 14'h3756: rddata <= 8'h0F; 14'h3757: rddata <= 8'h0F;
            14'h3758: rddata <= 8'hFF; 14'h3759: rddata <= 8'hFF; 14'h375A: rddata <= 8'hFF; 14'h375B: rddata <= 8'h0F;
            14'h375C: rddata <= 8'h0F; 14'h375D: rddata <= 8'h0F; 14'h375E: rddata <= 8'h0F; 14'h375F: rddata <= 8'h0F;
            14'h3760: rddata <= 8'h00; 14'h3761: rddata <= 8'h00; 14'h3762: rddata <= 8'h00; 14'h3763: rddata <= 8'hFF;
            14'h3764: rddata <= 8'hFF; 14'h3765: rddata <= 8'h0F; 14'h3766: rddata <= 8'h0F; 14'h3767: rddata <= 8'h0F;
            14'h3768: rddata <= 8'hF0; 14'h3769: rddata <= 8'hF0; 14'h376A: rddata <= 8'hF0; 14'h376B: rddata <= 8'hFF;
            14'h376C: rddata <= 8'hFF; 14'h376D: rddata <= 8'h0F; 14'h376E: rddata <= 8'h0F; 14'h376F: rddata <= 8'h0F;
            14'h3770: rddata <= 8'h0F; 14'h3771: rddata <= 8'h0F; 14'h3772: rddata <= 8'h0F; 14'h3773: rddata <= 8'hFF;
            14'h3774: rddata <= 8'hFF; 14'h3775: rddata <= 8'h0F; 14'h3776: rddata <= 8'h0F; 14'h3777: rddata <= 8'h0F;
            14'h3778: rddata <= 8'hFF; 14'h3779: rddata <= 8'hFF; 14'h377A: rddata <= 8'hFF; 14'h377B: rddata <= 8'hFF;
            14'h377C: rddata <= 8'hFF; 14'h377D: rddata <= 8'h0F; 14'h377E: rddata <= 8'h0F; 14'h377F: rddata <= 8'h0F;
            14'h3780: rddata <= 8'h00; 14'h3781: rddata <= 8'h00; 14'h3782: rddata <= 8'h00; 14'h3783: rddata <= 8'h00;
            14'h3784: rddata <= 8'h00; 14'h3785: rddata <= 8'hFF; 14'h3786: rddata <= 8'hFF; 14'h3787: rddata <= 8'hFF;
            14'h3788: rddata <= 8'hF0; 14'h3789: rddata <= 8'hF0; 14'h378A: rddata <= 8'hF0; 14'h378B: rddata <= 8'h00;
            14'h378C: rddata <= 8'h00; 14'h378D: rddata <= 8'hFF; 14'h378E: rddata <= 8'hFF; 14'h378F: rddata <= 8'hFF;
            14'h3790: rddata <= 8'h0F; 14'h3791: rddata <= 8'h0F; 14'h3792: rddata <= 8'h0F; 14'h3793: rddata <= 8'h00;
            14'h3794: rddata <= 8'h00; 14'h3795: rddata <= 8'hFF; 14'h3796: rddata <= 8'hFF; 14'h3797: rddata <= 8'hFF;
            14'h3798: rddata <= 8'hFF; 14'h3799: rddata <= 8'hFF; 14'h379A: rddata <= 8'hFF; 14'h379B: rddata <= 8'h00;
            14'h379C: rddata <= 8'h00; 14'h379D: rddata <= 8'hFF; 14'h379E: rddata <= 8'hFF; 14'h379F: rddata <= 8'hFF;
            14'h37A0: rddata <= 8'h00; 14'h37A1: rddata <= 8'h00; 14'h37A2: rddata <= 8'h00; 14'h37A3: rddata <= 8'hF0;
            14'h37A4: rddata <= 8'hF0; 14'h37A5: rddata <= 8'hFF; 14'h37A6: rddata <= 8'hFF; 14'h37A7: rddata <= 8'hFF;
            14'h37A8: rddata <= 8'hF0; 14'h37A9: rddata <= 8'hF0; 14'h37AA: rddata <= 8'hF0; 14'h37AB: rddata <= 8'hF0;
            14'h37AC: rddata <= 8'hF0; 14'h37AD: rddata <= 8'hFF; 14'h37AE: rddata <= 8'hFF; 14'h37AF: rddata <= 8'hFF;
            14'h37B0: rddata <= 8'h0F; 14'h37B1: rddata <= 8'h0F; 14'h37B2: rddata <= 8'h0F; 14'h37B3: rddata <= 8'hF0;
            14'h37B4: rddata <= 8'hF0; 14'h37B5: rddata <= 8'hFF; 14'h37B6: rddata <= 8'hFF; 14'h37B7: rddata <= 8'hFF;
            14'h37B8: rddata <= 8'hFF; 14'h37B9: rddata <= 8'hFF; 14'h37BA: rddata <= 8'hFF; 14'h37BB: rddata <= 8'hF0;
            14'h37BC: rddata <= 8'hF0; 14'h37BD: rddata <= 8'hFF; 14'h37BE: rddata <= 8'hFF; 14'h37BF: rddata <= 8'hFF;
            14'h37C0: rddata <= 8'h00; 14'h37C1: rddata <= 8'h00; 14'h37C2: rddata <= 8'h00; 14'h37C3: rddata <= 8'h0F;
            14'h37C4: rddata <= 8'h0F; 14'h37C5: rddata <= 8'hFF; 14'h37C6: rddata <= 8'hFF; 14'h37C7: rddata <= 8'hFF;
            14'h37C8: rddata <= 8'hF0; 14'h37C9: rddata <= 8'hF0; 14'h37CA: rddata <= 8'hF0; 14'h37CB: rddata <= 8'h0F;
            14'h37CC: rddata <= 8'h0F; 14'h37CD: rddata <= 8'hFF; 14'h37CE: rddata <= 8'hFF; 14'h37CF: rddata <= 8'hFF;
            14'h37D0: rddata <= 8'h0F; 14'h37D1: rddata <= 8'h0F; 14'h37D2: rddata <= 8'h0F; 14'h37D3: rddata <= 8'h0F;
            14'h37D4: rddata <= 8'h0F; 14'h37D5: rddata <= 8'hFF; 14'h37D6: rddata <= 8'hFF; 14'h37D7: rddata <= 8'hFF;
            14'h37D8: rddata <= 8'hFF; 14'h37D9: rddata <= 8'hFF; 14'h37DA: rddata <= 8'hFF; 14'h37DB: rddata <= 8'h0F;
            14'h37DC: rddata <= 8'h0F; 14'h37DD: rddata <= 8'hFF; 14'h37DE: rddata <= 8'hFF; 14'h37DF: rddata <= 8'hFF;
            14'h37E0: rddata <= 8'h00; 14'h37E1: rddata <= 8'h00; 14'h37E2: rddata <= 8'h00; 14'h37E3: rddata <= 8'hFF;
            14'h37E4: rddata <= 8'hFF; 14'h37E5: rddata <= 8'hFF; 14'h37E6: rddata <= 8'hFF; 14'h37E7: rddata <= 8'hFF;
            14'h37E8: rddata <= 8'hF0; 14'h37E9: rddata <= 8'hF0; 14'h37EA: rddata <= 8'hF0; 14'h37EB: rddata <= 8'hFF;
            14'h37EC: rddata <= 8'hFF; 14'h37ED: rddata <= 8'hFF; 14'h37EE: rddata <= 8'hFF; 14'h37EF: rddata <= 8'hFF;
            14'h37F0: rddata <= 8'h0F; 14'h37F1: rddata <= 8'h0F; 14'h37F2: rddata <= 8'h0F; 14'h37F3: rddata <= 8'hFF;
            14'h37F4: rddata <= 8'hFF; 14'h37F5: rddata <= 8'hFF; 14'h37F6: rddata <= 8'hFF; 14'h37F7: rddata <= 8'hFF;
            14'h37F8: rddata <= 8'hFF; 14'h37F9: rddata <= 8'hFF; 14'h37FA: rddata <= 8'hFF; 14'h37FB: rddata <= 8'hFF;
            14'h37FC: rddata <= 8'hFF; 14'h37FD: rddata <= 8'hFF; 14'h37FE: rddata <= 8'hFF; 14'h37FF: rddata <= 8'hFF;
            14'h3800: rddata <= 8'h00; 14'h3801: rddata <= 8'h00; 14'h3802: rddata <= 8'h00; 14'h3803: rddata <= 8'h00;
            14'h3804: rddata <= 8'h00; 14'h3805: rddata <= 8'h00; 14'h3806: rddata <= 8'h00; 14'h3807: rddata <= 8'h00;
            14'h3808: rddata <= 8'h7E; 14'h3809: rddata <= 8'h81; 14'h380A: rddata <= 8'hA5; 14'h380B: rddata <= 8'h81;
            14'h380C: rddata <= 8'hBD; 14'h380D: rddata <= 8'h99; 14'h380E: rddata <= 8'h81; 14'h380F: rddata <= 8'h7E;
            14'h3810: rddata <= 8'h7E; 14'h3811: rddata <= 8'hFF; 14'h3812: rddata <= 8'hDB; 14'h3813: rddata <= 8'hFF;
            14'h3814: rddata <= 8'hC3; 14'h3815: rddata <= 8'hE7; 14'h3816: rddata <= 8'hFF; 14'h3817: rddata <= 8'h7E;
            14'h3818: rddata <= 8'h36; 14'h3819: rddata <= 8'h7F; 14'h381A: rddata <= 8'h7F; 14'h381B: rddata <= 8'h7F;
            14'h381C: rddata <= 8'h3E; 14'h381D: rddata <= 8'h1C; 14'h381E: rddata <= 8'h08; 14'h381F: rddata <= 8'h00;
            14'h3820: rddata <= 8'h08; 14'h3821: rddata <= 8'h1C; 14'h3822: rddata <= 8'h3E; 14'h3823: rddata <= 8'h7F;
            14'h3824: rddata <= 8'h3E; 14'h3825: rddata <= 8'h1C; 14'h3826: rddata <= 8'h08; 14'h3827: rddata <= 8'h00;
            14'h3828: rddata <= 8'h18; 14'h3829: rddata <= 8'h3C; 14'h382A: rddata <= 8'h3C; 14'h382B: rddata <= 8'hE7;
            14'h382C: rddata <= 8'hE7; 14'h382D: rddata <= 8'hDB; 14'h382E: rddata <= 8'h18; 14'h382F: rddata <= 8'h3C;
            14'h3830: rddata <= 8'h18; 14'h3831: rddata <= 8'h3C; 14'h3832: rddata <= 8'h7E; 14'h3833: rddata <= 8'hFF;
            14'h3834: rddata <= 8'hFF; 14'h3835: rddata <= 8'hDB; 14'h3836: rddata <= 8'h18; 14'h3837: rddata <= 8'h3C;
            14'h3838: rddata <= 8'h00; 14'h3839: rddata <= 8'h00; 14'h383A: rddata <= 8'h18; 14'h383B: rddata <= 8'h3C;
            14'h383C: rddata <= 8'h3C; 14'h383D: rddata <= 8'h18; 14'h383E: rddata <= 8'h00; 14'h383F: rddata <= 8'h00;
            14'h3840: rddata <= 8'hFF; 14'h3841: rddata <= 8'hFF; 14'h3842: rddata <= 8'hE7; 14'h3843: rddata <= 8'hC3;
            14'h3844: rddata <= 8'hC3; 14'h3845: rddata <= 8'hE7; 14'h3846: rddata <= 8'hFF; 14'h3847: rddata <= 8'hFF;
            14'h3848: rddata <= 8'h00; 14'h3849: rddata <= 8'h3C; 14'h384A: rddata <= 8'h66; 14'h384B: rddata <= 8'h42;
            14'h384C: rddata <= 8'h42; 14'h384D: rddata <= 8'h66; 14'h384E: rddata <= 8'h3C; 14'h384F: rddata <= 8'h00;
            14'h3850: rddata <= 8'hFF; 14'h3851: rddata <= 8'hC3; 14'h3852: rddata <= 8'h99; 14'h3853: rddata <= 8'hBD;
            14'h3854: rddata <= 8'hBD; 14'h3855: rddata <= 8'h99; 14'h3856: rddata <= 8'hC3; 14'h3857: rddata <= 8'hFF;
            14'h3858: rddata <= 8'h0F; 14'h3859: rddata <= 8'h07; 14'h385A: rddata <= 8'h0F; 14'h385B: rddata <= 8'h7D;
            14'h385C: rddata <= 8'hCC; 14'h385D: rddata <= 8'hCC; 14'h385E: rddata <= 8'hCC; 14'h385F: rddata <= 8'h78;
            14'h3860: rddata <= 8'h3C; 14'h3861: rddata <= 8'h66; 14'h3862: rddata <= 8'h66; 14'h3863: rddata <= 8'h66;
            14'h3864: rddata <= 8'h3C; 14'h3865: rddata <= 8'h18; 14'h3866: rddata <= 8'h7E; 14'h3867: rddata <= 8'h18;
            14'h3868: rddata <= 8'h3F; 14'h3869: rddata <= 8'h33; 14'h386A: rddata <= 8'h3F; 14'h386B: rddata <= 8'h30;
            14'h386C: rddata <= 8'h30; 14'h386D: rddata <= 8'h70; 14'h386E: rddata <= 8'hF0; 14'h386F: rddata <= 8'hE0;
            14'h3870: rddata <= 8'h7F; 14'h3871: rddata <= 8'h63; 14'h3872: rddata <= 8'h7F; 14'h3873: rddata <= 8'h63;
            14'h3874: rddata <= 8'h63; 14'h3875: rddata <= 8'h67; 14'h3876: rddata <= 8'hE6; 14'h3877: rddata <= 8'hC0;
            14'h3878: rddata <= 8'h99; 14'h3879: rddata <= 8'h5A; 14'h387A: rddata <= 8'h3C; 14'h387B: rddata <= 8'hE7;
            14'h387C: rddata <= 8'hE7; 14'h387D: rddata <= 8'h3C; 14'h387E: rddata <= 8'h5A; 14'h387F: rddata <= 8'h99;
            14'h3880: rddata <= 8'h80; 14'h3881: rddata <= 8'hE0; 14'h3882: rddata <= 8'hF8; 14'h3883: rddata <= 8'hFE;
            14'h3884: rddata <= 8'hF8; 14'h3885: rddata <= 8'hE0; 14'h3886: rddata <= 8'h80; 14'h3887: rddata <= 8'h00;
            14'h3888: rddata <= 8'h02; 14'h3889: rddata <= 8'h0E; 14'h388A: rddata <= 8'h3E; 14'h388B: rddata <= 8'hFE;
            14'h388C: rddata <= 8'h3E; 14'h388D: rddata <= 8'h0E; 14'h388E: rddata <= 8'h02; 14'h388F: rddata <= 8'h00;
            14'h3890: rddata <= 8'h18; 14'h3891: rddata <= 8'h3C; 14'h3892: rddata <= 8'h7E; 14'h3893: rddata <= 8'h18;
            14'h3894: rddata <= 8'h18; 14'h3895: rddata <= 8'h7E; 14'h3896: rddata <= 8'h3C; 14'h3897: rddata <= 8'h18;
            14'h3898: rddata <= 8'h66; 14'h3899: rddata <= 8'h66; 14'h389A: rddata <= 8'h66; 14'h389B: rddata <= 8'h66;
            14'h389C: rddata <= 8'h66; 14'h389D: rddata <= 8'h00; 14'h389E: rddata <= 8'h66; 14'h389F: rddata <= 8'h00;
            14'h38A0: rddata <= 8'h7F; 14'h38A1: rddata <= 8'hDB; 14'h38A2: rddata <= 8'hDB; 14'h38A3: rddata <= 8'h7B;
            14'h38A4: rddata <= 8'h1B; 14'h38A5: rddata <= 8'h1B; 14'h38A6: rddata <= 8'h1B; 14'h38A7: rddata <= 8'h00;
            14'h38A8: rddata <= 8'h3C; 14'h38A9: rddata <= 8'h66; 14'h38AA: rddata <= 8'h38; 14'h38AB: rddata <= 8'h6C;
            14'h38AC: rddata <= 8'h6C; 14'h38AD: rddata <= 8'h38; 14'h38AE: rddata <= 8'hCC; 14'h38AF: rddata <= 8'h78;
            14'h38B0: rddata <= 8'h00; 14'h38B1: rddata <= 8'h00; 14'h38B2: rddata <= 8'h00; 14'h38B3: rddata <= 8'h00;
            14'h38B4: rddata <= 8'h7E; 14'h38B5: rddata <= 8'h7E; 14'h38B6: rddata <= 8'h7E; 14'h38B7: rddata <= 8'h00;
            14'h38B8: rddata <= 8'h18; 14'h38B9: rddata <= 8'h3C; 14'h38BA: rddata <= 8'h7E; 14'h38BB: rddata <= 8'h18;
            14'h38BC: rddata <= 8'h7E; 14'h38BD: rddata <= 8'h3C; 14'h38BE: rddata <= 8'h18; 14'h38BF: rddata <= 8'hFF;
            14'h38C0: rddata <= 8'h18; 14'h38C1: rddata <= 8'h3C; 14'h38C2: rddata <= 8'h7E; 14'h38C3: rddata <= 8'h18;
            14'h38C4: rddata <= 8'h18; 14'h38C5: rddata <= 8'h18; 14'h38C6: rddata <= 8'h18; 14'h38C7: rddata <= 8'h00;
            14'h38C8: rddata <= 8'h18; 14'h38C9: rddata <= 8'h18; 14'h38CA: rddata <= 8'h18; 14'h38CB: rddata <= 8'h18;
            14'h38CC: rddata <= 8'h7E; 14'h38CD: rddata <= 8'h3C; 14'h38CE: rddata <= 8'h18; 14'h38CF: rddata <= 8'h00;
            14'h38D0: rddata <= 8'h00; 14'h38D1: rddata <= 8'h08; 14'h38D2: rddata <= 8'h0C; 14'h38D3: rddata <= 8'hFE;
            14'h38D4: rddata <= 8'hFE; 14'h38D5: rddata <= 8'h0C; 14'h38D6: rddata <= 8'h08; 14'h38D7: rddata <= 8'h00;
            14'h38D8: rddata <= 8'h00; 14'h38D9: rddata <= 8'h10; 14'h38DA: rddata <= 8'h30; 14'h38DB: rddata <= 8'h7F;
            14'h38DC: rddata <= 8'h7F; 14'h38DD: rddata <= 8'h30; 14'h38DE: rddata <= 8'h10; 14'h38DF: rddata <= 8'h00;
            14'h38E0: rddata <= 8'h00; 14'h38E1: rddata <= 8'h00; 14'h38E2: rddata <= 8'hC0; 14'h38E3: rddata <= 8'hC0;
            14'h38E4: rddata <= 8'hC0; 14'h38E5: rddata <= 8'hFE; 14'h38E6: rddata <= 8'h00; 14'h38E7: rddata <= 8'h00;
            14'h38E8: rddata <= 8'h00; 14'h38E9: rddata <= 8'h24; 14'h38EA: rddata <= 8'h66; 14'h38EB: rddata <= 8'hFF;
            14'h38EC: rddata <= 8'h66; 14'h38ED: rddata <= 8'h24; 14'h38EE: rddata <= 8'h00; 14'h38EF: rddata <= 8'h00;
            14'h38F0: rddata <= 8'h00; 14'h38F1: rddata <= 8'h18; 14'h38F2: rddata <= 8'h3C; 14'h38F3: rddata <= 8'h7E;
            14'h38F4: rddata <= 8'hFF; 14'h38F5: rddata <= 8'hFF; 14'h38F6: rddata <= 8'h00; 14'h38F7: rddata <= 8'h00;
            14'h38F8: rddata <= 8'h00; 14'h38F9: rddata <= 8'hFF; 14'h38FA: rddata <= 8'hFF; 14'h38FB: rddata <= 8'h7E;
            14'h38FC: rddata <= 8'h3C; 14'h38FD: rddata <= 8'h18; 14'h38FE: rddata <= 8'h00; 14'h38FF: rddata <= 8'h00;
            14'h3900: rddata <= 8'h00; 14'h3901: rddata <= 8'h00; 14'h3902: rddata <= 8'h00; 14'h3903: rddata <= 8'h00;
            14'h3904: rddata <= 8'h00; 14'h3905: rddata <= 8'h00; 14'h3906: rddata <= 8'h00; 14'h3907: rddata <= 8'h00;
            14'h3908: rddata <= 8'h18; 14'h3909: rddata <= 8'h18; 14'h390A: rddata <= 8'h18; 14'h390B: rddata <= 8'h18;
            14'h390C: rddata <= 8'h00; 14'h390D: rddata <= 8'h00; 14'h390E: rddata <= 8'h18; 14'h390F: rddata <= 8'h00;
            14'h3910: rddata <= 8'h66; 14'h3911: rddata <= 8'h66; 14'h3912: rddata <= 8'h66; 14'h3913: rddata <= 8'h00;
            14'h3914: rddata <= 8'h00; 14'h3915: rddata <= 8'h00; 14'h3916: rddata <= 8'h00; 14'h3917: rddata <= 8'h00;
            14'h3918: rddata <= 8'h6C; 14'h3919: rddata <= 8'h6C; 14'h391A: rddata <= 8'hFE; 14'h391B: rddata <= 8'h6C;
            14'h391C: rddata <= 8'hFE; 14'h391D: rddata <= 8'h6C; 14'h391E: rddata <= 8'h6C; 14'h391F: rddata <= 8'h00;
            14'h3920: rddata <= 8'h18; 14'h3921: rddata <= 8'h3E; 14'h3922: rddata <= 8'h60; 14'h3923: rddata <= 8'h3C;
            14'h3924: rddata <= 8'h06; 14'h3925: rddata <= 8'h7C; 14'h3926: rddata <= 8'h18; 14'h3927: rddata <= 8'h00;
            14'h3928: rddata <= 8'h62; 14'h3929: rddata <= 8'h66; 14'h392A: rddata <= 8'h0C; 14'h392B: rddata <= 8'h18;
            14'h392C: rddata <= 8'h30; 14'h392D: rddata <= 8'h66; 14'h392E: rddata <= 8'h46; 14'h392F: rddata <= 8'h00;
            14'h3930: rddata <= 8'h38; 14'h3931: rddata <= 8'h6C; 14'h3932: rddata <= 8'h38; 14'h3933: rddata <= 8'h76;
            14'h3934: rddata <= 8'hDC; 14'h3935: rddata <= 8'hCC; 14'h3936: rddata <= 8'h76; 14'h3937: rddata <= 8'h00;
            14'h3938: rddata <= 8'h18; 14'h3939: rddata <= 8'h18; 14'h393A: rddata <= 8'h30; 14'h393B: rddata <= 8'h00;
            14'h393C: rddata <= 8'h00; 14'h393D: rddata <= 8'h00; 14'h393E: rddata <= 8'h00; 14'h393F: rddata <= 8'h00;
            14'h3940: rddata <= 8'h0C; 14'h3941: rddata <= 8'h18; 14'h3942: rddata <= 8'h30; 14'h3943: rddata <= 8'h30;
            14'h3944: rddata <= 8'h30; 14'h3945: rddata <= 8'h18; 14'h3946: rddata <= 8'h0C; 14'h3947: rddata <= 8'h00;
            14'h3948: rddata <= 8'h30; 14'h3949: rddata <= 8'h18; 14'h394A: rddata <= 8'h0C; 14'h394B: rddata <= 8'h0C;
            14'h394C: rddata <= 8'h0C; 14'h394D: rddata <= 8'h18; 14'h394E: rddata <= 8'h30; 14'h394F: rddata <= 8'h00;
            14'h3950: rddata <= 8'h00; 14'h3951: rddata <= 8'h66; 14'h3952: rddata <= 8'h3C; 14'h3953: rddata <= 8'hFF;
            14'h3954: rddata <= 8'h3C; 14'h3955: rddata <= 8'h66; 14'h3956: rddata <= 8'h00; 14'h3957: rddata <= 8'h00;
            14'h3958: rddata <= 8'h00; 14'h3959: rddata <= 8'h18; 14'h395A: rddata <= 8'h18; 14'h395B: rddata <= 8'h7E;
            14'h395C: rddata <= 8'h18; 14'h395D: rddata <= 8'h18; 14'h395E: rddata <= 8'h00; 14'h395F: rddata <= 8'h00;
            14'h3960: rddata <= 8'h00; 14'h3961: rddata <= 8'h00; 14'h3962: rddata <= 8'h00; 14'h3963: rddata <= 8'h00;
            14'h3964: rddata <= 8'h00; 14'h3965: rddata <= 8'h18; 14'h3966: rddata <= 8'h18; 14'h3967: rddata <= 8'h30;
            14'h3968: rddata <= 8'h00; 14'h3969: rddata <= 8'h00; 14'h396A: rddata <= 8'h00; 14'h396B: rddata <= 8'h7E;
            14'h396C: rddata <= 8'h00; 14'h396D: rddata <= 8'h00; 14'h396E: rddata <= 8'h00; 14'h396F: rddata <= 8'h00;
            14'h3970: rddata <= 8'h00; 14'h3971: rddata <= 8'h00; 14'h3972: rddata <= 8'h00; 14'h3973: rddata <= 8'h00;
            14'h3974: rddata <= 8'h00; 14'h3975: rddata <= 8'h18; 14'h3976: rddata <= 8'h18; 14'h3977: rddata <= 8'h00;
            14'h3978: rddata <= 8'h06; 14'h3979: rddata <= 8'h0C; 14'h397A: rddata <= 8'h18; 14'h397B: rddata <= 8'h30;
            14'h397C: rddata <= 8'h60; 14'h397D: rddata <= 8'hC0; 14'h397E: rddata <= 8'h80; 14'h397F: rddata <= 8'h00;
            14'h3980: rddata <= 8'h3C; 14'h3981: rddata <= 8'h66; 14'h3982: rddata <= 8'h6E; 14'h3983: rddata <= 8'h76;
            14'h3984: rddata <= 8'h66; 14'h3985: rddata <= 8'h66; 14'h3986: rddata <= 8'h3C; 14'h3987: rddata <= 8'h00;
            14'h3988: rddata <= 8'h18; 14'h3989: rddata <= 8'h18; 14'h398A: rddata <= 8'h38; 14'h398B: rddata <= 8'h18;
            14'h398C: rddata <= 8'h18; 14'h398D: rddata <= 8'h18; 14'h398E: rddata <= 8'h7E; 14'h398F: rddata <= 8'h00;
            14'h3990: rddata <= 8'h3C; 14'h3991: rddata <= 8'h66; 14'h3992: rddata <= 8'h06; 14'h3993: rddata <= 8'h0C;
            14'h3994: rddata <= 8'h30; 14'h3995: rddata <= 8'h60; 14'h3996: rddata <= 8'h7E; 14'h3997: rddata <= 8'h00;
            14'h3998: rddata <= 8'h3C; 14'h3999: rddata <= 8'h66; 14'h399A: rddata <= 8'h06; 14'h399B: rddata <= 8'h1C;
            14'h399C: rddata <= 8'h06; 14'h399D: rddata <= 8'h66; 14'h399E: rddata <= 8'h3C; 14'h399F: rddata <= 8'h00;
            14'h39A0: rddata <= 8'h0E; 14'h39A1: rddata <= 8'h1E; 14'h39A2: rddata <= 8'h36; 14'h39A3: rddata <= 8'h66;
            14'h39A4: rddata <= 8'h7F; 14'h39A5: rddata <= 8'h06; 14'h39A6: rddata <= 8'h06; 14'h39A7: rddata <= 8'h00;
            14'h39A8: rddata <= 8'h7E; 14'h39A9: rddata <= 8'h60; 14'h39AA: rddata <= 8'h7C; 14'h39AB: rddata <= 8'h06;
            14'h39AC: rddata <= 8'h06; 14'h39AD: rddata <= 8'h66; 14'h39AE: rddata <= 8'h3C; 14'h39AF: rddata <= 8'h00;
            14'h39B0: rddata <= 8'h3C; 14'h39B1: rddata <= 8'h66; 14'h39B2: rddata <= 8'h60; 14'h39B3: rddata <= 8'h7C;
            14'h39B4: rddata <= 8'h66; 14'h39B5: rddata <= 8'h66; 14'h39B6: rddata <= 8'h3C; 14'h39B7: rddata <= 8'h00;
            14'h39B8: rddata <= 8'h7E; 14'h39B9: rddata <= 8'h66; 14'h39BA: rddata <= 8'h06; 14'h39BB: rddata <= 8'h0C;
            14'h39BC: rddata <= 8'h18; 14'h39BD: rddata <= 8'h18; 14'h39BE: rddata <= 8'h18; 14'h39BF: rddata <= 8'h00;
            14'h39C0: rddata <= 8'h3C; 14'h39C1: rddata <= 8'h66; 14'h39C2: rddata <= 8'h66; 14'h39C3: rddata <= 8'h3C;
            14'h39C4: rddata <= 8'h66; 14'h39C5: rddata <= 8'h66; 14'h39C6: rddata <= 8'h3C; 14'h39C7: rddata <= 8'h00;
            14'h39C8: rddata <= 8'h3C; 14'h39C9: rddata <= 8'h66; 14'h39CA: rddata <= 8'h66; 14'h39CB: rddata <= 8'h3E;
            14'h39CC: rddata <= 8'h06; 14'h39CD: rddata <= 8'h66; 14'h39CE: rddata <= 8'h3C; 14'h39CF: rddata <= 8'h00;
            14'h39D0: rddata <= 8'h00; 14'h39D1: rddata <= 8'h18; 14'h39D2: rddata <= 8'h18; 14'h39D3: rddata <= 8'h00;
            14'h39D4: rddata <= 8'h00; 14'h39D5: rddata <= 8'h18; 14'h39D6: rddata <= 8'h18; 14'h39D7: rddata <= 8'h00;
            14'h39D8: rddata <= 8'h00; 14'h39D9: rddata <= 8'h18; 14'h39DA: rddata <= 8'h18; 14'h39DB: rddata <= 8'h00;
            14'h39DC: rddata <= 8'h00; 14'h39DD: rddata <= 8'h18; 14'h39DE: rddata <= 8'h18; 14'h39DF: rddata <= 8'h30;
            14'h39E0: rddata <= 8'h0C; 14'h39E1: rddata <= 8'h18; 14'h39E2: rddata <= 8'h30; 14'h39E3: rddata <= 8'h60;
            14'h39E4: rddata <= 8'h30; 14'h39E5: rddata <= 8'h18; 14'h39E6: rddata <= 8'h0C; 14'h39E7: rddata <= 8'h00;
            14'h39E8: rddata <= 8'h00; 14'h39E9: rddata <= 8'h00; 14'h39EA: rddata <= 8'h7E; 14'h39EB: rddata <= 8'h00;
            14'h39EC: rddata <= 8'h7E; 14'h39ED: rddata <= 8'h00; 14'h39EE: rddata <= 8'h00; 14'h39EF: rddata <= 8'h00;
            14'h39F0: rddata <= 8'h30; 14'h39F1: rddata <= 8'h18; 14'h39F2: rddata <= 8'h0C; 14'h39F3: rddata <= 8'h06;
            14'h39F4: rddata <= 8'h0C; 14'h39F5: rddata <= 8'h18; 14'h39F6: rddata <= 8'h30; 14'h39F7: rddata <= 8'h00;
            14'h39F8: rddata <= 8'h3C; 14'h39F9: rddata <= 8'h66; 14'h39FA: rddata <= 8'h06; 14'h39FB: rddata <= 8'h0C;
            14'h39FC: rddata <= 8'h18; 14'h39FD: rddata <= 8'h00; 14'h39FE: rddata <= 8'h18; 14'h39FF: rddata <= 8'h00;
            14'h3A00: rddata <= 8'h3C; 14'h3A01: rddata <= 8'h66; 14'h3A02: rddata <= 8'h6E; 14'h3A03: rddata <= 8'h6E;
            14'h3A04: rddata <= 8'h60; 14'h3A05: rddata <= 8'h62; 14'h3A06: rddata <= 8'h3C; 14'h3A07: rddata <= 8'h00;
            14'h3A08: rddata <= 8'h18; 14'h3A09: rddata <= 8'h3C; 14'h3A0A: rddata <= 8'h66; 14'h3A0B: rddata <= 8'h7E;
            14'h3A0C: rddata <= 8'h66; 14'h3A0D: rddata <= 8'h66; 14'h3A0E: rddata <= 8'h66; 14'h3A0F: rddata <= 8'h00;
            14'h3A10: rddata <= 8'h7C; 14'h3A11: rddata <= 8'h66; 14'h3A12: rddata <= 8'h66; 14'h3A13: rddata <= 8'h7C;
            14'h3A14: rddata <= 8'h66; 14'h3A15: rddata <= 8'h66; 14'h3A16: rddata <= 8'h7C; 14'h3A17: rddata <= 8'h00;
            14'h3A18: rddata <= 8'h3C; 14'h3A19: rddata <= 8'h66; 14'h3A1A: rddata <= 8'h60; 14'h3A1B: rddata <= 8'h60;
            14'h3A1C: rddata <= 8'h60; 14'h3A1D: rddata <= 8'h66; 14'h3A1E: rddata <= 8'h3C; 14'h3A1F: rddata <= 8'h00;
            14'h3A20: rddata <= 8'h78; 14'h3A21: rddata <= 8'h6C; 14'h3A22: rddata <= 8'h66; 14'h3A23: rddata <= 8'h66;
            14'h3A24: rddata <= 8'h66; 14'h3A25: rddata <= 8'h6C; 14'h3A26: rddata <= 8'h78; 14'h3A27: rddata <= 8'h00;
            14'h3A28: rddata <= 8'h7E; 14'h3A29: rddata <= 8'h60; 14'h3A2A: rddata <= 8'h60; 14'h3A2B: rddata <= 8'h78;
            14'h3A2C: rddata <= 8'h60; 14'h3A2D: rddata <= 8'h60; 14'h3A2E: rddata <= 8'h7E; 14'h3A2F: rddata <= 8'h00;
            14'h3A30: rddata <= 8'h7E; 14'h3A31: rddata <= 8'h60; 14'h3A32: rddata <= 8'h60; 14'h3A33: rddata <= 8'h78;
            14'h3A34: rddata <= 8'h60; 14'h3A35: rddata <= 8'h60; 14'h3A36: rddata <= 8'h60; 14'h3A37: rddata <= 8'h00;
            14'h3A38: rddata <= 8'h3C; 14'h3A39: rddata <= 8'h66; 14'h3A3A: rddata <= 8'h60; 14'h3A3B: rddata <= 8'h6E;
            14'h3A3C: rddata <= 8'h66; 14'h3A3D: rddata <= 8'h66; 14'h3A3E: rddata <= 8'h3C; 14'h3A3F: rddata <= 8'h00;
            14'h3A40: rddata <= 8'h66; 14'h3A41: rddata <= 8'h66; 14'h3A42: rddata <= 8'h66; 14'h3A43: rddata <= 8'h7E;
            14'h3A44: rddata <= 8'h66; 14'h3A45: rddata <= 8'h66; 14'h3A46: rddata <= 8'h66; 14'h3A47: rddata <= 8'h00;
            14'h3A48: rddata <= 8'h3C; 14'h3A49: rddata <= 8'h18; 14'h3A4A: rddata <= 8'h18; 14'h3A4B: rddata <= 8'h18;
            14'h3A4C: rddata <= 8'h18; 14'h3A4D: rddata <= 8'h18; 14'h3A4E: rddata <= 8'h3C; 14'h3A4F: rddata <= 8'h00;
            14'h3A50: rddata <= 8'h1E; 14'h3A51: rddata <= 8'h0C; 14'h3A52: rddata <= 8'h0C; 14'h3A53: rddata <= 8'h0C;
            14'h3A54: rddata <= 8'h0C; 14'h3A55: rddata <= 8'h6C; 14'h3A56: rddata <= 8'h38; 14'h3A57: rddata <= 8'h00;
            14'h3A58: rddata <= 8'h66; 14'h3A59: rddata <= 8'h6C; 14'h3A5A: rddata <= 8'h78; 14'h3A5B: rddata <= 8'h70;
            14'h3A5C: rddata <= 8'h78; 14'h3A5D: rddata <= 8'h6C; 14'h3A5E: rddata <= 8'h66; 14'h3A5F: rddata <= 8'h00;
            14'h3A60: rddata <= 8'h60; 14'h3A61: rddata <= 8'h60; 14'h3A62: rddata <= 8'h60; 14'h3A63: rddata <= 8'h60;
            14'h3A64: rddata <= 8'h60; 14'h3A65: rddata <= 8'h60; 14'h3A66: rddata <= 8'h7E; 14'h3A67: rddata <= 8'h00;
            14'h3A68: rddata <= 8'h63; 14'h3A69: rddata <= 8'h77; 14'h3A6A: rddata <= 8'h7F; 14'h3A6B: rddata <= 8'h6B;
            14'h3A6C: rddata <= 8'h63; 14'h3A6D: rddata <= 8'h63; 14'h3A6E: rddata <= 8'h63; 14'h3A6F: rddata <= 8'h00;
            14'h3A70: rddata <= 8'h66; 14'h3A71: rddata <= 8'h76; 14'h3A72: rddata <= 8'h7E; 14'h3A73: rddata <= 8'h7E;
            14'h3A74: rddata <= 8'h6E; 14'h3A75: rddata <= 8'h66; 14'h3A76: rddata <= 8'h66; 14'h3A77: rddata <= 8'h00;
            14'h3A78: rddata <= 8'h3C; 14'h3A79: rddata <= 8'h66; 14'h3A7A: rddata <= 8'h66; 14'h3A7B: rddata <= 8'h66;
            14'h3A7C: rddata <= 8'h66; 14'h3A7D: rddata <= 8'h66; 14'h3A7E: rddata <= 8'h3C; 14'h3A7F: rddata <= 8'h00;
            14'h3A80: rddata <= 8'h7C; 14'h3A81: rddata <= 8'h66; 14'h3A82: rddata <= 8'h66; 14'h3A83: rddata <= 8'h7C;
            14'h3A84: rddata <= 8'h60; 14'h3A85: rddata <= 8'h60; 14'h3A86: rddata <= 8'h60; 14'h3A87: rddata <= 8'h00;
            14'h3A88: rddata <= 8'h3C; 14'h3A89: rddata <= 8'h66; 14'h3A8A: rddata <= 8'h66; 14'h3A8B: rddata <= 8'h66;
            14'h3A8C: rddata <= 8'h66; 14'h3A8D: rddata <= 8'h3C; 14'h3A8E: rddata <= 8'h0E; 14'h3A8F: rddata <= 8'h00;
            14'h3A90: rddata <= 8'h7C; 14'h3A91: rddata <= 8'h66; 14'h3A92: rddata <= 8'h66; 14'h3A93: rddata <= 8'h7C;
            14'h3A94: rddata <= 8'h78; 14'h3A95: rddata <= 8'h6C; 14'h3A96: rddata <= 8'h66; 14'h3A97: rddata <= 8'h00;
            14'h3A98: rddata <= 8'h3C; 14'h3A99: rddata <= 8'h66; 14'h3A9A: rddata <= 8'h60; 14'h3A9B: rddata <= 8'h3C;
            14'h3A9C: rddata <= 8'h06; 14'h3A9D: rddata <= 8'h66; 14'h3A9E: rddata <= 8'h3C; 14'h3A9F: rddata <= 8'h00;
            14'h3AA0: rddata <= 8'h7E; 14'h3AA1: rddata <= 8'h18; 14'h3AA2: rddata <= 8'h18; 14'h3AA3: rddata <= 8'h18;
            14'h3AA4: rddata <= 8'h18; 14'h3AA5: rddata <= 8'h18; 14'h3AA6: rddata <= 8'h18; 14'h3AA7: rddata <= 8'h00;
            14'h3AA8: rddata <= 8'h66; 14'h3AA9: rddata <= 8'h66; 14'h3AAA: rddata <= 8'h66; 14'h3AAB: rddata <= 8'h66;
            14'h3AAC: rddata <= 8'h66; 14'h3AAD: rddata <= 8'h66; 14'h3AAE: rddata <= 8'h3C; 14'h3AAF: rddata <= 8'h00;
            14'h3AB0: rddata <= 8'h66; 14'h3AB1: rddata <= 8'h66; 14'h3AB2: rddata <= 8'h66; 14'h3AB3: rddata <= 8'h66;
            14'h3AB4: rddata <= 8'h66; 14'h3AB5: rddata <= 8'h3C; 14'h3AB6: rddata <= 8'h18; 14'h3AB7: rddata <= 8'h00;
            14'h3AB8: rddata <= 8'h63; 14'h3AB9: rddata <= 8'h63; 14'h3ABA: rddata <= 8'h63; 14'h3ABB: rddata <= 8'h6B;
            14'h3ABC: rddata <= 8'h7F; 14'h3ABD: rddata <= 8'h77; 14'h3ABE: rddata <= 8'h63; 14'h3ABF: rddata <= 8'h00;
            14'h3AC0: rddata <= 8'h66; 14'h3AC1: rddata <= 8'h66; 14'h3AC2: rddata <= 8'h3C; 14'h3AC3: rddata <= 8'h18;
            14'h3AC4: rddata <= 8'h3C; 14'h3AC5: rddata <= 8'h66; 14'h3AC6: rddata <= 8'h66; 14'h3AC7: rddata <= 8'h00;
            14'h3AC8: rddata <= 8'h66; 14'h3AC9: rddata <= 8'h66; 14'h3ACA: rddata <= 8'h66; 14'h3ACB: rddata <= 8'h3C;
            14'h3ACC: rddata <= 8'h18; 14'h3ACD: rddata <= 8'h18; 14'h3ACE: rddata <= 8'h18; 14'h3ACF: rddata <= 8'h00;
            14'h3AD0: rddata <= 8'h7E; 14'h3AD1: rddata <= 8'h06; 14'h3AD2: rddata <= 8'h0C; 14'h3AD3: rddata <= 8'h18;
            14'h3AD4: rddata <= 8'h30; 14'h3AD5: rddata <= 8'h60; 14'h3AD6: rddata <= 8'h7E; 14'h3AD7: rddata <= 8'h00;
            14'h3AD8: rddata <= 8'h3C; 14'h3AD9: rddata <= 8'h30; 14'h3ADA: rddata <= 8'h30; 14'h3ADB: rddata <= 8'h30;
            14'h3ADC: rddata <= 8'h30; 14'h3ADD: rddata <= 8'h30; 14'h3ADE: rddata <= 8'h3C; 14'h3ADF: rddata <= 8'h00;
            14'h3AE0: rddata <= 8'hC0; 14'h3AE1: rddata <= 8'h60; 14'h3AE2: rddata <= 8'h30; 14'h3AE3: rddata <= 8'h18;
            14'h3AE4: rddata <= 8'h0C; 14'h3AE5: rddata <= 8'h06; 14'h3AE6: rddata <= 8'h02; 14'h3AE7: rddata <= 8'h00;
            14'h3AE8: rddata <= 8'h3C; 14'h3AE9: rddata <= 8'h0C; 14'h3AEA: rddata <= 8'h0C; 14'h3AEB: rddata <= 8'h0C;
            14'h3AEC: rddata <= 8'h0C; 14'h3AED: rddata <= 8'h0C; 14'h3AEE: rddata <= 8'h3C; 14'h3AEF: rddata <= 8'h00;
            14'h3AF0: rddata <= 8'h10; 14'h3AF1: rddata <= 8'h38; 14'h3AF2: rddata <= 8'h6C; 14'h3AF3: rddata <= 8'hC6;
            14'h3AF4: rddata <= 8'h00; 14'h3AF5: rddata <= 8'h00; 14'h3AF6: rddata <= 8'h00; 14'h3AF7: rddata <= 8'h00;
            14'h3AF8: rddata <= 8'h00; 14'h3AF9: rddata <= 8'h00; 14'h3AFA: rddata <= 8'h00; 14'h3AFB: rddata <= 8'h00;
            14'h3AFC: rddata <= 8'h00; 14'h3AFD: rddata <= 8'h00; 14'h3AFE: rddata <= 8'hFE; 14'h3AFF: rddata <= 8'h00;
            14'h3B00: rddata <= 8'h30; 14'h3B01: rddata <= 8'h30; 14'h3B02: rddata <= 8'h18; 14'h3B03: rddata <= 8'h00;
            14'h3B04: rddata <= 8'h00; 14'h3B05: rddata <= 8'h00; 14'h3B06: rddata <= 8'h00; 14'h3B07: rddata <= 8'h00;
            14'h3B08: rddata <= 8'h00; 14'h3B09: rddata <= 8'h00; 14'h3B0A: rddata <= 8'h3C; 14'h3B0B: rddata <= 8'h06;
            14'h3B0C: rddata <= 8'h3E; 14'h3B0D: rddata <= 8'h66; 14'h3B0E: rddata <= 8'h3E; 14'h3B0F: rddata <= 8'h00;
            14'h3B10: rddata <= 8'h60; 14'h3B11: rddata <= 8'h60; 14'h3B12: rddata <= 8'h7C; 14'h3B13: rddata <= 8'h66;
            14'h3B14: rddata <= 8'h66; 14'h3B15: rddata <= 8'h66; 14'h3B16: rddata <= 8'h7C; 14'h3B17: rddata <= 8'h00;
            14'h3B18: rddata <= 8'h00; 14'h3B19: rddata <= 8'h00; 14'h3B1A: rddata <= 8'h3C; 14'h3B1B: rddata <= 8'h60;
            14'h3B1C: rddata <= 8'h60; 14'h3B1D: rddata <= 8'h60; 14'h3B1E: rddata <= 8'h3C; 14'h3B1F: rddata <= 8'h00;
            14'h3B20: rddata <= 8'h06; 14'h3B21: rddata <= 8'h06; 14'h3B22: rddata <= 8'h3E; 14'h3B23: rddata <= 8'h66;
            14'h3B24: rddata <= 8'h66; 14'h3B25: rddata <= 8'h66; 14'h3B26: rddata <= 8'h3E; 14'h3B27: rddata <= 8'h00;
            14'h3B28: rddata <= 8'h00; 14'h3B29: rddata <= 8'h00; 14'h3B2A: rddata <= 8'h3C; 14'h3B2B: rddata <= 8'h66;
            14'h3B2C: rddata <= 8'h7E; 14'h3B2D: rddata <= 8'h60; 14'h3B2E: rddata <= 8'h3C; 14'h3B2F: rddata <= 8'h00;
            14'h3B30: rddata <= 8'h0E; 14'h3B31: rddata <= 8'h18; 14'h3B32: rddata <= 8'h18; 14'h3B33: rddata <= 8'h3E;
            14'h3B34: rddata <= 8'h18; 14'h3B35: rddata <= 8'h18; 14'h3B36: rddata <= 8'h18; 14'h3B37: rddata <= 8'h00;
            14'h3B38: rddata <= 8'h00; 14'h3B39: rddata <= 8'h00; 14'h3B3A: rddata <= 8'h3E; 14'h3B3B: rddata <= 8'h66;
            14'h3B3C: rddata <= 8'h66; 14'h3B3D: rddata <= 8'h3E; 14'h3B3E: rddata <= 8'h06; 14'h3B3F: rddata <= 8'h7C;
            14'h3B40: rddata <= 8'h60; 14'h3B41: rddata <= 8'h60; 14'h3B42: rddata <= 8'h7C; 14'h3B43: rddata <= 8'h66;
            14'h3B44: rddata <= 8'h66; 14'h3B45: rddata <= 8'h66; 14'h3B46: rddata <= 8'h66; 14'h3B47: rddata <= 8'h00;
            14'h3B48: rddata <= 8'h18; 14'h3B49: rddata <= 8'h00; 14'h3B4A: rddata <= 8'h38; 14'h3B4B: rddata <= 8'h18;
            14'h3B4C: rddata <= 8'h18; 14'h3B4D: rddata <= 8'h18; 14'h3B4E: rddata <= 8'h3C; 14'h3B4F: rddata <= 8'h00;
            14'h3B50: rddata <= 8'h18; 14'h3B51: rddata <= 8'h00; 14'h3B52: rddata <= 8'h38; 14'h3B53: rddata <= 8'h18;
            14'h3B54: rddata <= 8'h18; 14'h3B55: rddata <= 8'h18; 14'h3B56: rddata <= 8'h18; 14'h3B57: rddata <= 8'h70;
            14'h3B58: rddata <= 8'h60; 14'h3B59: rddata <= 8'h60; 14'h3B5A: rddata <= 8'h66; 14'h3B5B: rddata <= 8'h6C;
            14'h3B5C: rddata <= 8'h78; 14'h3B5D: rddata <= 8'h6C; 14'h3B5E: rddata <= 8'h66; 14'h3B5F: rddata <= 8'h00;
            14'h3B60: rddata <= 8'h38; 14'h3B61: rddata <= 8'h18; 14'h3B62: rddata <= 8'h18; 14'h3B63: rddata <= 8'h18;
            14'h3B64: rddata <= 8'h18; 14'h3B65: rddata <= 8'h18; 14'h3B66: rddata <= 8'h3C; 14'h3B67: rddata <= 8'h00;
            14'h3B68: rddata <= 8'h00; 14'h3B69: rddata <= 8'h00; 14'h3B6A: rddata <= 8'h66; 14'h3B6B: rddata <= 8'h7F;
            14'h3B6C: rddata <= 8'h7F; 14'h3B6D: rddata <= 8'h6B; 14'h3B6E: rddata <= 8'h63; 14'h3B6F: rddata <= 8'h00;
            14'h3B70: rddata <= 8'h00; 14'h3B71: rddata <= 8'h00; 14'h3B72: rddata <= 8'h7C; 14'h3B73: rddata <= 8'h66;
            14'h3B74: rddata <= 8'h66; 14'h3B75: rddata <= 8'h66; 14'h3B76: rddata <= 8'h66; 14'h3B77: rddata <= 8'h00;
            14'h3B78: rddata <= 8'h00; 14'h3B79: rddata <= 8'h00; 14'h3B7A: rddata <= 8'h3C; 14'h3B7B: rddata <= 8'h66;
            14'h3B7C: rddata <= 8'h66; 14'h3B7D: rddata <= 8'h66; 14'h3B7E: rddata <= 8'h3C; 14'h3B7F: rddata <= 8'h00;
            14'h3B80: rddata <= 8'h00; 14'h3B81: rddata <= 8'h00; 14'h3B82: rddata <= 8'h7C; 14'h3B83: rddata <= 8'h66;
            14'h3B84: rddata <= 8'h66; 14'h3B85: rddata <= 8'h7C; 14'h3B86: rddata <= 8'h60; 14'h3B87: rddata <= 8'h60;
            14'h3B88: rddata <= 8'h00; 14'h3B89: rddata <= 8'h00; 14'h3B8A: rddata <= 8'h3E; 14'h3B8B: rddata <= 8'h66;
            14'h3B8C: rddata <= 8'h66; 14'h3B8D: rddata <= 8'h3E; 14'h3B8E: rddata <= 8'h06; 14'h3B8F: rddata <= 8'h06;
            14'h3B90: rddata <= 8'h00; 14'h3B91: rddata <= 8'h00; 14'h3B92: rddata <= 8'h7C; 14'h3B93: rddata <= 8'h66;
            14'h3B94: rddata <= 8'h60; 14'h3B95: rddata <= 8'h60; 14'h3B96: rddata <= 8'h60; 14'h3B97: rddata <= 8'h00;
            14'h3B98: rddata <= 8'h00; 14'h3B99: rddata <= 8'h00; 14'h3B9A: rddata <= 8'h3E; 14'h3B9B: rddata <= 8'h60;
            14'h3B9C: rddata <= 8'h3C; 14'h3B9D: rddata <= 8'h06; 14'h3B9E: rddata <= 8'h7C; 14'h3B9F: rddata <= 8'h00;
            14'h3BA0: rddata <= 8'h18; 14'h3BA1: rddata <= 8'h18; 14'h3BA2: rddata <= 8'h7E; 14'h3BA3: rddata <= 8'h18;
            14'h3BA4: rddata <= 8'h18; 14'h3BA5: rddata <= 8'h18; 14'h3BA6: rddata <= 8'h0E; 14'h3BA7: rddata <= 8'h00;
            14'h3BA8: rddata <= 8'h00; 14'h3BA9: rddata <= 8'h00; 14'h3BAA: rddata <= 8'h66; 14'h3BAB: rddata <= 8'h66;
            14'h3BAC: rddata <= 8'h66; 14'h3BAD: rddata <= 8'h66; 14'h3BAE: rddata <= 8'h3E; 14'h3BAF: rddata <= 8'h00;
            14'h3BB0: rddata <= 8'h00; 14'h3BB1: rddata <= 8'h00; 14'h3BB2: rddata <= 8'h66; 14'h3BB3: rddata <= 8'h66;
            14'h3BB4: rddata <= 8'h66; 14'h3BB5: rddata <= 8'h3C; 14'h3BB6: rddata <= 8'h18; 14'h3BB7: rddata <= 8'h00;
            14'h3BB8: rddata <= 8'h00; 14'h3BB9: rddata <= 8'h00; 14'h3BBA: rddata <= 8'h63; 14'h3BBB: rddata <= 8'h6B;
            14'h3BBC: rddata <= 8'h7F; 14'h3BBD: rddata <= 8'h3E; 14'h3BBE: rddata <= 8'h36; 14'h3BBF: rddata <= 8'h00;
            14'h3BC0: rddata <= 8'h00; 14'h3BC1: rddata <= 8'h00; 14'h3BC2: rddata <= 8'h66; 14'h3BC3: rddata <= 8'h3C;
            14'h3BC4: rddata <= 8'h18; 14'h3BC5: rddata <= 8'h3C; 14'h3BC6: rddata <= 8'h66; 14'h3BC7: rddata <= 8'h00;
            14'h3BC8: rddata <= 8'h00; 14'h3BC9: rddata <= 8'h00; 14'h3BCA: rddata <= 8'h66; 14'h3BCB: rddata <= 8'h66;
            14'h3BCC: rddata <= 8'h66; 14'h3BCD: rddata <= 8'h3E; 14'h3BCE: rddata <= 8'h0C; 14'h3BCF: rddata <= 8'h78;
            14'h3BD0: rddata <= 8'h00; 14'h3BD1: rddata <= 8'h00; 14'h3BD2: rddata <= 8'h7E; 14'h3BD3: rddata <= 8'h0C;
            14'h3BD4: rddata <= 8'h18; 14'h3BD5: rddata <= 8'h30; 14'h3BD6: rddata <= 8'h7E; 14'h3BD7: rddata <= 8'h00;
            14'h3BD8: rddata <= 8'h0E; 14'h3BD9: rddata <= 8'h18; 14'h3BDA: rddata <= 8'h18; 14'h3BDB: rddata <= 8'h70;
            14'h3BDC: rddata <= 8'h18; 14'h3BDD: rddata <= 8'h18; 14'h3BDE: rddata <= 8'h0E; 14'h3BDF: rddata <= 8'h00;
            14'h3BE0: rddata <= 8'h18; 14'h3BE1: rddata <= 8'h18; 14'h3BE2: rddata <= 8'h18; 14'h3BE3: rddata <= 8'h00;
            14'h3BE4: rddata <= 8'h18; 14'h3BE5: rddata <= 8'h18; 14'h3BE6: rddata <= 8'h18; 14'h3BE7: rddata <= 8'h00;
            14'h3BE8: rddata <= 8'h70; 14'h3BE9: rddata <= 8'h18; 14'h3BEA: rddata <= 8'h18; 14'h3BEB: rddata <= 8'h0E;
            14'h3BEC: rddata <= 8'h18; 14'h3BED: rddata <= 8'h18; 14'h3BEE: rddata <= 8'h70; 14'h3BEF: rddata <= 8'h00;
            14'h3BF0: rddata <= 8'h00; 14'h3BF1: rddata <= 8'h00; 14'h3BF2: rddata <= 8'h76; 14'h3BF3: rddata <= 8'hDC;
            14'h3BF4: rddata <= 8'h00; 14'h3BF5: rddata <= 8'h00; 14'h3BF6: rddata <= 8'h00; 14'h3BF7: rddata <= 8'h00;
            14'h3BF8: rddata <= 8'h00; 14'h3BF9: rddata <= 8'h10; 14'h3BFA: rddata <= 8'h38; 14'h3BFB: rddata <= 8'h6C;
            14'h3BFC: rddata <= 8'hC6; 14'h3BFD: rddata <= 8'hC6; 14'h3BFE: rddata <= 8'hFE; 14'h3BFF: rddata <= 8'h00;
            14'h3C00: rddata <= 8'h78; 14'h3C01: rddata <= 8'hCC; 14'h3C02: rddata <= 8'hC0; 14'h3C03: rddata <= 8'hCC;
            14'h3C04: rddata <= 8'h78; 14'h3C05: rddata <= 8'h18; 14'h3C06: rddata <= 8'h0C; 14'h3C07: rddata <= 8'h78;
            14'h3C08: rddata <= 8'h00; 14'h3C09: rddata <= 8'h66; 14'h3C0A: rddata <= 8'h00; 14'h3C0B: rddata <= 8'h66;
            14'h3C0C: rddata <= 8'h66; 14'h3C0D: rddata <= 8'h66; 14'h3C0E: rddata <= 8'h3E; 14'h3C0F: rddata <= 8'h00;
            14'h3C10: rddata <= 8'h0E; 14'h3C11: rddata <= 8'h00; 14'h3C12: rddata <= 8'h3C; 14'h3C13: rddata <= 8'h66;
            14'h3C14: rddata <= 8'h7E; 14'h3C15: rddata <= 8'h60; 14'h3C16: rddata <= 8'h3C; 14'h3C17: rddata <= 8'h00;
            14'h3C18: rddata <= 8'h3C; 14'h3C19: rddata <= 8'h42; 14'h3C1A: rddata <= 8'h3C; 14'h3C1B: rddata <= 8'h06;
            14'h3C1C: rddata <= 8'h3E; 14'h3C1D: rddata <= 8'h66; 14'h3C1E: rddata <= 8'h3E; 14'h3C1F: rddata <= 8'h00;
            14'h3C20: rddata <= 8'h66; 14'h3C21: rddata <= 8'h00; 14'h3C22: rddata <= 8'h3C; 14'h3C23: rddata <= 8'h06;
            14'h3C24: rddata <= 8'h3E; 14'h3C25: rddata <= 8'h66; 14'h3C26: rddata <= 8'h3E; 14'h3C27: rddata <= 8'h00;
            14'h3C28: rddata <= 8'h70; 14'h3C29: rddata <= 8'h00; 14'h3C2A: rddata <= 8'h3C; 14'h3C2B: rddata <= 8'h06;
            14'h3C2C: rddata <= 8'h3E; 14'h3C2D: rddata <= 8'h66; 14'h3C2E: rddata <= 8'h3E; 14'h3C2F: rddata <= 8'h00;
            14'h3C30: rddata <= 8'h18; 14'h3C31: rddata <= 8'h18; 14'h3C32: rddata <= 8'h3C; 14'h3C33: rddata <= 8'h06;
            14'h3C34: rddata <= 8'h3E; 14'h3C35: rddata <= 8'h66; 14'h3C36: rddata <= 8'h3E; 14'h3C37: rddata <= 8'h00;
            14'h3C38: rddata <= 8'h00; 14'h3C39: rddata <= 8'h00; 14'h3C3A: rddata <= 8'h3C; 14'h3C3B: rddata <= 8'h60;
            14'h3C3C: rddata <= 8'h60; 14'h3C3D: rddata <= 8'h3C; 14'h3C3E: rddata <= 8'h06; 14'h3C3F: rddata <= 8'h1C;
            14'h3C40: rddata <= 8'h7E; 14'h3C41: rddata <= 8'hC3; 14'h3C42: rddata <= 8'h3C; 14'h3C43: rddata <= 8'h66;
            14'h3C44: rddata <= 8'h7E; 14'h3C45: rddata <= 8'h60; 14'h3C46: rddata <= 8'h3C; 14'h3C47: rddata <= 8'h00;
            14'h3C48: rddata <= 8'h66; 14'h3C49: rddata <= 8'h00; 14'h3C4A: rddata <= 8'h3C; 14'h3C4B: rddata <= 8'h66;
            14'h3C4C: rddata <= 8'h7E; 14'h3C4D: rddata <= 8'h60; 14'h3C4E: rddata <= 8'h3C; 14'h3C4F: rddata <= 8'h00;
            14'h3C50: rddata <= 8'h70; 14'h3C51: rddata <= 8'h00; 14'h3C52: rddata <= 8'h3C; 14'h3C53: rddata <= 8'h66;
            14'h3C54: rddata <= 8'h7E; 14'h3C55: rddata <= 8'h60; 14'h3C56: rddata <= 8'h3C; 14'h3C57: rddata <= 8'h00;
            14'h3C58: rddata <= 8'h00; 14'h3C59: rddata <= 8'h66; 14'h3C5A: rddata <= 8'h00; 14'h3C5B: rddata <= 8'h38;
            14'h3C5C: rddata <= 8'h18; 14'h3C5D: rddata <= 8'h18; 14'h3C5E: rddata <= 8'h3C; 14'h3C5F: rddata <= 8'h00;
            14'h3C60: rddata <= 8'h18; 14'h3C61: rddata <= 8'h24; 14'h3C62: rddata <= 8'h00; 14'h3C63: rddata <= 8'h38;
            14'h3C64: rddata <= 8'h18; 14'h3C65: rddata <= 8'h18; 14'h3C66: rddata <= 8'h3C; 14'h3C67: rddata <= 8'h00;
            14'h3C68: rddata <= 8'h20; 14'h3C69: rddata <= 8'h10; 14'h3C6A: rddata <= 8'h00; 14'h3C6B: rddata <= 8'h38;
            14'h3C6C: rddata <= 8'h18; 14'h3C6D: rddata <= 8'h18; 14'h3C6E: rddata <= 8'h3C; 14'h3C6F: rddata <= 8'h00;
            14'h3C70: rddata <= 8'h5A; 14'h3C71: rddata <= 8'h3C; 14'h3C72: rddata <= 8'h66; 14'h3C73: rddata <= 8'h7E;
            14'h3C74: rddata <= 8'h66; 14'h3C75: rddata <= 8'h66; 14'h3C76: rddata <= 8'h66; 14'h3C77: rddata <= 8'h00;
            14'h3C78: rddata <= 8'h18; 14'h3C79: rddata <= 8'h18; 14'h3C7A: rddata <= 8'h00; 14'h3C7B: rddata <= 8'h3C;
            14'h3C7C: rddata <= 8'h66; 14'h3C7D: rddata <= 8'h7E; 14'h3C7E: rddata <= 8'h66; 14'h3C7F: rddata <= 8'h00;
            14'h3C80: rddata <= 8'h1C; 14'h3C81: rddata <= 8'h00; 14'h3C82: rddata <= 8'h7E; 14'h3C83: rddata <= 8'h60;
            14'h3C84: rddata <= 8'h78; 14'h3C85: rddata <= 8'h60; 14'h3C86: rddata <= 8'h7E; 14'h3C87: rddata <= 8'h00;
            14'h3C88: rddata <= 8'h00; 14'h3C89: rddata <= 8'h00; 14'h3C8A: rddata <= 8'h7F; 14'h3C8B: rddata <= 8'h0C;
            14'h3C8C: rddata <= 8'h7F; 14'h3C8D: rddata <= 8'hCC; 14'h3C8E: rddata <= 8'h7F; 14'h3C8F: rddata <= 8'h00;
            14'h3C90: rddata <= 8'h3E; 14'h3C91: rddata <= 8'h6C; 14'h3C92: rddata <= 8'hCC; 14'h3C93: rddata <= 8'hFE;
            14'h3C94: rddata <= 8'hCC; 14'h3C95: rddata <= 8'hCC; 14'h3C96: rddata <= 8'hCE; 14'h3C97: rddata <= 8'h00;
            14'h3C98: rddata <= 8'h3C; 14'h3C99: rddata <= 8'h66; 14'h3C9A: rddata <= 8'h00; 14'h3C9B: rddata <= 8'h3C;
            14'h3C9C: rddata <= 8'h66; 14'h3C9D: rddata <= 8'h66; 14'h3C9E: rddata <= 8'h3C; 14'h3C9F: rddata <= 8'h00;
            14'h3CA0: rddata <= 8'h00; 14'h3CA1: rddata <= 8'h66; 14'h3CA2: rddata <= 8'h00; 14'h3CA3: rddata <= 8'h3C;
            14'h3CA4: rddata <= 8'h66; 14'h3CA5: rddata <= 8'h66; 14'h3CA6: rddata <= 8'h3C; 14'h3CA7: rddata <= 8'h00;
            14'h3CA8: rddata <= 8'h00; 14'h3CA9: rddata <= 8'h70; 14'h3CAA: rddata <= 8'h00; 14'h3CAB: rddata <= 8'h3C;
            14'h3CAC: rddata <= 8'h66; 14'h3CAD: rddata <= 8'h66; 14'h3CAE: rddata <= 8'h3C; 14'h3CAF: rddata <= 8'h00;
            14'h3CB0: rddata <= 8'h3C; 14'h3CB1: rddata <= 8'h66; 14'h3CB2: rddata <= 8'h00; 14'h3CB3: rddata <= 8'h66;
            14'h3CB4: rddata <= 8'h66; 14'h3CB5: rddata <= 8'h66; 14'h3CB6: rddata <= 8'h3E; 14'h3CB7: rddata <= 8'h00;
            14'h3CB8: rddata <= 8'h00; 14'h3CB9: rddata <= 8'h70; 14'h3CBA: rddata <= 8'h00; 14'h3CBB: rddata <= 8'h66;
            14'h3CBC: rddata <= 8'h66; 14'h3CBD: rddata <= 8'h66; 14'h3CBE: rddata <= 8'h3E; 14'h3CBF: rddata <= 8'h00;
            14'h3CC0: rddata <= 8'h00; 14'h3CC1: rddata <= 8'h66; 14'h3CC2: rddata <= 8'h00; 14'h3CC3: rddata <= 8'h66;
            14'h3CC4: rddata <= 8'h66; 14'h3CC5: rddata <= 8'h3E; 14'h3CC6: rddata <= 8'h0C; 14'h3CC7: rddata <= 8'h78;
            14'h3CC8: rddata <= 8'hC3; 14'h3CC9: rddata <= 8'h3C; 14'h3CCA: rddata <= 8'h66; 14'h3CCB: rddata <= 8'h66;
            14'h3CCC: rddata <= 8'h66; 14'h3CCD: rddata <= 8'h66; 14'h3CCE: rddata <= 8'h3C; 14'h3CCF: rddata <= 8'h00;
            14'h3CD0: rddata <= 8'h66; 14'h3CD1: rddata <= 8'h00; 14'h3CD2: rddata <= 8'h66; 14'h3CD3: rddata <= 8'h66;
            14'h3CD4: rddata <= 8'h66; 14'h3CD5: rddata <= 8'h66; 14'h3CD6: rddata <= 8'h3C; 14'h3CD7: rddata <= 8'h00;
            14'h3CD8: rddata <= 8'h18; 14'h3CD9: rddata <= 8'h18; 14'h3CDA: rddata <= 8'h7E; 14'h3CDB: rddata <= 8'hC0;
            14'h3CDC: rddata <= 8'hC0; 14'h3CDD: rddata <= 8'h7E; 14'h3CDE: rddata <= 8'h18; 14'h3CDF: rddata <= 8'h18;
            14'h3CE0: rddata <= 8'h0C; 14'h3CE1: rddata <= 8'h12; 14'h3CE2: rddata <= 8'h30; 14'h3CE3: rddata <= 8'h7C;
            14'h3CE4: rddata <= 8'h30; 14'h3CE5: rddata <= 8'h62; 14'h3CE6: rddata <= 8'hFC; 14'h3CE7: rddata <= 8'h00;
            14'h3CE8: rddata <= 8'hCC; 14'h3CE9: rddata <= 8'hCC; 14'h3CEA: rddata <= 8'h78; 14'h3CEB: rddata <= 8'hFC;
            14'h3CEC: rddata <= 8'h30; 14'h3CED: rddata <= 8'hFC; 14'h3CEE: rddata <= 8'h30; 14'h3CEF: rddata <= 8'h30;
            14'h3CF0: rddata <= 8'hF8; 14'h3CF1: rddata <= 8'hCC; 14'h3CF2: rddata <= 8'hCC; 14'h3CF3: rddata <= 8'hFA;
            14'h3CF4: rddata <= 8'hC6; 14'h3CF5: rddata <= 8'hCF; 14'h3CF6: rddata <= 8'hC6; 14'h3CF7: rddata <= 8'hC7;
            14'h3CF8: rddata <= 8'h0E; 14'h3CF9: rddata <= 8'h1B; 14'h3CFA: rddata <= 8'h18; 14'h3CFB: rddata <= 8'h3C;
            14'h3CFC: rddata <= 8'h18; 14'h3CFD: rddata <= 8'h18; 14'h3CFE: rddata <= 8'hD8; 14'h3CFF: rddata <= 8'h70;
            14'h3D00: rddata <= 8'h0E; 14'h3D01: rddata <= 8'h00; 14'h3D02: rddata <= 8'h3C; 14'h3D03: rddata <= 8'h06;
            14'h3D04: rddata <= 8'h3E; 14'h3D05: rddata <= 8'h66; 14'h3D06: rddata <= 8'h3E; 14'h3D07: rddata <= 8'h00;
            14'h3D08: rddata <= 8'h08; 14'h3D09: rddata <= 8'h10; 14'h3D0A: rddata <= 8'h00; 14'h3D0B: rddata <= 8'h38;
            14'h3D0C: rddata <= 8'h18; 14'h3D0D: rddata <= 8'h18; 14'h3D0E: rddata <= 8'h3C; 14'h3D0F: rddata <= 8'h00;
            14'h3D10: rddata <= 8'h00; 14'h3D11: rddata <= 8'h0E; 14'h3D12: rddata <= 8'h00; 14'h3D13: rddata <= 8'h3C;
            14'h3D14: rddata <= 8'h66; 14'h3D15: rddata <= 8'h66; 14'h3D16: rddata <= 8'h3C; 14'h3D17: rddata <= 8'h00;
            14'h3D18: rddata <= 8'h00; 14'h3D19: rddata <= 8'h0E; 14'h3D1A: rddata <= 8'h00; 14'h3D1B: rddata <= 8'h66;
            14'h3D1C: rddata <= 8'h66; 14'h3D1D: rddata <= 8'h66; 14'h3D1E: rddata <= 8'h3E; 14'h3D1F: rddata <= 8'h00;
            14'h3D20: rddata <= 8'h00; 14'h3D21: rddata <= 8'h7C; 14'h3D22: rddata <= 8'h00; 14'h3D23: rddata <= 8'h7C;
            14'h3D24: rddata <= 8'h66; 14'h3D25: rddata <= 8'h66; 14'h3D26: rddata <= 8'h66; 14'h3D27: rddata <= 8'h00;
            14'h3D28: rddata <= 8'h7E; 14'h3D29: rddata <= 8'h00; 14'h3D2A: rddata <= 8'h66; 14'h3D2B: rddata <= 8'h76;
            14'h3D2C: rddata <= 8'h7E; 14'h3D2D: rddata <= 8'h6E; 14'h3D2E: rddata <= 8'h66; 14'h3D2F: rddata <= 8'h00;
            14'h3D30: rddata <= 8'h3C; 14'h3D31: rddata <= 8'h6C; 14'h3D32: rddata <= 8'h6C; 14'h3D33: rddata <= 8'h3E;
            14'h3D34: rddata <= 8'h00; 14'h3D35: rddata <= 8'h7E; 14'h3D36: rddata <= 8'h00; 14'h3D37: rddata <= 8'h00;
            14'h3D38: rddata <= 8'h38; 14'h3D39: rddata <= 8'h6C; 14'h3D3A: rddata <= 8'h6C; 14'h3D3B: rddata <= 8'h38;
            14'h3D3C: rddata <= 8'h00; 14'h3D3D: rddata <= 8'h7C; 14'h3D3E: rddata <= 8'h00; 14'h3D3F: rddata <= 8'h00;
            14'h3D40: rddata <= 8'h18; 14'h3D41: rddata <= 8'h00; 14'h3D42: rddata <= 8'h18; 14'h3D43: rddata <= 8'h30;
            14'h3D44: rddata <= 8'h60; 14'h3D45: rddata <= 8'h66; 14'h3D46: rddata <= 8'h3C; 14'h3D47: rddata <= 8'h00;
            14'h3D48: rddata <= 8'h00; 14'h3D49: rddata <= 8'h00; 14'h3D4A: rddata <= 8'h00; 14'h3D4B: rddata <= 8'h7E;
            14'h3D4C: rddata <= 8'h60; 14'h3D4D: rddata <= 8'h60; 14'h3D4E: rddata <= 8'h00; 14'h3D4F: rddata <= 8'h00;
            14'h3D50: rddata <= 8'h00; 14'h3D51: rddata <= 8'h00; 14'h3D52: rddata <= 8'h00; 14'h3D53: rddata <= 8'h7E;
            14'h3D54: rddata <= 8'h06; 14'h3D55: rddata <= 8'h06; 14'h3D56: rddata <= 8'h00; 14'h3D57: rddata <= 8'h00;
            14'h3D58: rddata <= 8'hC3; 14'h3D59: rddata <= 8'hC6; 14'h3D5A: rddata <= 8'hCC; 14'h3D5B: rddata <= 8'hDE;
            14'h3D5C: rddata <= 8'h33; 14'h3D5D: rddata <= 8'h66; 14'h3D5E: rddata <= 8'hCC; 14'h3D5F: rddata <= 8'h0F;
            14'h3D60: rddata <= 8'hC3; 14'h3D61: rddata <= 8'hC6; 14'h3D62: rddata <= 8'hCC; 14'h3D63: rddata <= 8'hDB;
            14'h3D64: rddata <= 8'h37; 14'h3D65: rddata <= 8'h6F; 14'h3D66: rddata <= 8'hCF; 14'h3D67: rddata <= 8'h03;
            14'h3D68: rddata <= 8'h18; 14'h3D69: rddata <= 8'h18; 14'h3D6A: rddata <= 8'h00; 14'h3D6B: rddata <= 8'h18;
            14'h3D6C: rddata <= 8'h18; 14'h3D6D: rddata <= 8'h18; 14'h3D6E: rddata <= 8'h18; 14'h3D6F: rddata <= 8'h00;
            14'h3D70: rddata <= 8'h00; 14'h3D71: rddata <= 8'h33; 14'h3D72: rddata <= 8'h66; 14'h3D73: rddata <= 8'hCC;
            14'h3D74: rddata <= 8'h66; 14'h3D75: rddata <= 8'h33; 14'h3D76: rddata <= 8'h00; 14'h3D77: rddata <= 8'h00;
            14'h3D78: rddata <= 8'h00; 14'h3D79: rddata <= 8'hCC; 14'h3D7A: rddata <= 8'h66; 14'h3D7B: rddata <= 8'h33;
            14'h3D7C: rddata <= 8'h66; 14'h3D7D: rddata <= 8'hCC; 14'h3D7E: rddata <= 8'h00; 14'h3D7F: rddata <= 8'h00;
            14'h3D80: rddata <= 8'h22; 14'h3D81: rddata <= 8'h88; 14'h3D82: rddata <= 8'h22; 14'h3D83: rddata <= 8'h88;
            14'h3D84: rddata <= 8'h22; 14'h3D85: rddata <= 8'h88; 14'h3D86: rddata <= 8'h22; 14'h3D87: rddata <= 8'h88;
            14'h3D88: rddata <= 8'h55; 14'h3D89: rddata <= 8'hAA; 14'h3D8A: rddata <= 8'h55; 14'h3D8B: rddata <= 8'hAA;
            14'h3D8C: rddata <= 8'h55; 14'h3D8D: rddata <= 8'hAA; 14'h3D8E: rddata <= 8'h55; 14'h3D8F: rddata <= 8'hAA;
            14'h3D90: rddata <= 8'hBB; 14'h3D91: rddata <= 8'hEE; 14'h3D92: rddata <= 8'hBB; 14'h3D93: rddata <= 8'hEE;
            14'h3D94: rddata <= 8'hBB; 14'h3D95: rddata <= 8'hEE; 14'h3D96: rddata <= 8'hBB; 14'h3D97: rddata <= 8'hEE;
            14'h3D98: rddata <= 8'h18; 14'h3D99: rddata <= 8'h18; 14'h3D9A: rddata <= 8'h18; 14'h3D9B: rddata <= 8'h18;
            14'h3D9C: rddata <= 8'h18; 14'h3D9D: rddata <= 8'h18; 14'h3D9E: rddata <= 8'h18; 14'h3D9F: rddata <= 8'h18;
            14'h3DA0: rddata <= 8'h18; 14'h3DA1: rddata <= 8'h18; 14'h3DA2: rddata <= 8'h18; 14'h3DA3: rddata <= 8'h18;
            14'h3DA4: rddata <= 8'hF8; 14'h3DA5: rddata <= 8'h18; 14'h3DA6: rddata <= 8'h18; 14'h3DA7: rddata <= 8'h18;
            14'h3DA8: rddata <= 8'h18; 14'h3DA9: rddata <= 8'h18; 14'h3DAA: rddata <= 8'hF8; 14'h3DAB: rddata <= 8'h18;
            14'h3DAC: rddata <= 8'hF8; 14'h3DAD: rddata <= 8'h18; 14'h3DAE: rddata <= 8'h18; 14'h3DAF: rddata <= 8'h18;
            14'h3DB0: rddata <= 8'h36; 14'h3DB1: rddata <= 8'h36; 14'h3DB2: rddata <= 8'h36; 14'h3DB3: rddata <= 8'h36;
            14'h3DB4: rddata <= 8'hF6; 14'h3DB5: rddata <= 8'h36; 14'h3DB6: rddata <= 8'h36; 14'h3DB7: rddata <= 8'h36;
            14'h3DB8: rddata <= 8'h00; 14'h3DB9: rddata <= 8'h00; 14'h3DBA: rddata <= 8'h00; 14'h3DBB: rddata <= 8'h00;
            14'h3DBC: rddata <= 8'hFE; 14'h3DBD: rddata <= 8'h36; 14'h3DBE: rddata <= 8'h36; 14'h3DBF: rddata <= 8'h36;
            14'h3DC0: rddata <= 8'h00; 14'h3DC1: rddata <= 8'h00; 14'h3DC2: rddata <= 8'hF8; 14'h3DC3: rddata <= 8'h18;
            14'h3DC4: rddata <= 8'hF8; 14'h3DC5: rddata <= 8'h18; 14'h3DC6: rddata <= 8'h18; 14'h3DC7: rddata <= 8'h18;
            14'h3DC8: rddata <= 8'h36; 14'h3DC9: rddata <= 8'h36; 14'h3DCA: rddata <= 8'hF6; 14'h3DCB: rddata <= 8'h06;
            14'h3DCC: rddata <= 8'hF6; 14'h3DCD: rddata <= 8'h36; 14'h3DCE: rddata <= 8'h36; 14'h3DCF: rddata <= 8'h36;
            14'h3DD0: rddata <= 8'h36; 14'h3DD1: rddata <= 8'h36; 14'h3DD2: rddata <= 8'h36; 14'h3DD3: rddata <= 8'h36;
            14'h3DD4: rddata <= 8'h36; 14'h3DD5: rddata <= 8'h36; 14'h3DD6: rddata <= 8'h36; 14'h3DD7: rddata <= 8'h36;
            14'h3DD8: rddata <= 8'h00; 14'h3DD9: rddata <= 8'h00; 14'h3DDA: rddata <= 8'hFE; 14'h3DDB: rddata <= 8'h06;
            14'h3DDC: rddata <= 8'hF6; 14'h3DDD: rddata <= 8'h36; 14'h3DDE: rddata <= 8'h36; 14'h3DDF: rddata <= 8'h36;
            14'h3DE0: rddata <= 8'h36; 14'h3DE1: rddata <= 8'h36; 14'h3DE2: rddata <= 8'hF6; 14'h3DE3: rddata <= 8'h06;
            14'h3DE4: rddata <= 8'hFE; 14'h3DE5: rddata <= 8'h00; 14'h3DE6: rddata <= 8'h00; 14'h3DE7: rddata <= 8'h00;
            14'h3DE8: rddata <= 8'h36; 14'h3DE9: rddata <= 8'h36; 14'h3DEA: rddata <= 8'h36; 14'h3DEB: rddata <= 8'h36;
            14'h3DEC: rddata <= 8'hFE; 14'h3DED: rddata <= 8'h00; 14'h3DEE: rddata <= 8'h00; 14'h3DEF: rddata <= 8'h00;
            14'h3DF0: rddata <= 8'h18; 14'h3DF1: rddata <= 8'h18; 14'h3DF2: rddata <= 8'hF8; 14'h3DF3: rddata <= 8'h18;
            14'h3DF4: rddata <= 8'hF8; 14'h3DF5: rddata <= 8'h00; 14'h3DF6: rddata <= 8'h00; 14'h3DF7: rddata <= 8'h00;
            14'h3DF8: rddata <= 8'h00; 14'h3DF9: rddata <= 8'h00; 14'h3DFA: rddata <= 8'h00; 14'h3DFB: rddata <= 8'h00;
            14'h3DFC: rddata <= 8'hF8; 14'h3DFD: rddata <= 8'h18; 14'h3DFE: rddata <= 8'h18; 14'h3DFF: rddata <= 8'h18;
            14'h3E00: rddata <= 8'h18; 14'h3E01: rddata <= 8'h18; 14'h3E02: rddata <= 8'h18; 14'h3E03: rddata <= 8'h18;
            14'h3E04: rddata <= 8'h1F; 14'h3E05: rddata <= 8'h00; 14'h3E06: rddata <= 8'h00; 14'h3E07: rddata <= 8'h00;
            14'h3E08: rddata <= 8'h18; 14'h3E09: rddata <= 8'h18; 14'h3E0A: rddata <= 8'h18; 14'h3E0B: rddata <= 8'h18;
            14'h3E0C: rddata <= 8'hFF; 14'h3E0D: rddata <= 8'h00; 14'h3E0E: rddata <= 8'h00; 14'h3E0F: rddata <= 8'h00;
            14'h3E10: rddata <= 8'h00; 14'h3E11: rddata <= 8'h00; 14'h3E12: rddata <= 8'h00; 14'h3E13: rddata <= 8'h00;
            14'h3E14: rddata <= 8'hFF; 14'h3E15: rddata <= 8'h18; 14'h3E16: rddata <= 8'h18; 14'h3E17: rddata <= 8'h18;
            14'h3E18: rddata <= 8'h18; 14'h3E19: rddata <= 8'h18; 14'h3E1A: rddata <= 8'h18; 14'h3E1B: rddata <= 8'h18;
            14'h3E1C: rddata <= 8'h1F; 14'h3E1D: rddata <= 8'h18; 14'h3E1E: rddata <= 8'h18; 14'h3E1F: rddata <= 8'h18;
            14'h3E20: rddata <= 8'h00; 14'h3E21: rddata <= 8'h00; 14'h3E22: rddata <= 8'h00; 14'h3E23: rddata <= 8'h00;
            14'h3E24: rddata <= 8'hFF; 14'h3E25: rddata <= 8'h00; 14'h3E26: rddata <= 8'h00; 14'h3E27: rddata <= 8'h00;
            14'h3E28: rddata <= 8'h18; 14'h3E29: rddata <= 8'h18; 14'h3E2A: rddata <= 8'h18; 14'h3E2B: rddata <= 8'h18;
            14'h3E2C: rddata <= 8'hFF; 14'h3E2D: rddata <= 8'h18; 14'h3E2E: rddata <= 8'h18; 14'h3E2F: rddata <= 8'h18;
            14'h3E30: rddata <= 8'h18; 14'h3E31: rddata <= 8'h18; 14'h3E32: rddata <= 8'h1F; 14'h3E33: rddata <= 8'h18;
            14'h3E34: rddata <= 8'h1F; 14'h3E35: rddata <= 8'h18; 14'h3E36: rddata <= 8'h18; 14'h3E37: rddata <= 8'h18;
            14'h3E38: rddata <= 8'h36; 14'h3E39: rddata <= 8'h36; 14'h3E3A: rddata <= 8'h36; 14'h3E3B: rddata <= 8'h36;
            14'h3E3C: rddata <= 8'h37; 14'h3E3D: rddata <= 8'h36; 14'h3E3E: rddata <= 8'h36; 14'h3E3F: rddata <= 8'h36;
            14'h3E40: rddata <= 8'h36; 14'h3E41: rddata <= 8'h36; 14'h3E42: rddata <= 8'h37; 14'h3E43: rddata <= 8'h30;
            14'h3E44: rddata <= 8'h3F; 14'h3E45: rddata <= 8'h00; 14'h3E46: rddata <= 8'h00; 14'h3E47: rddata <= 8'h00;
            14'h3E48: rddata <= 8'h00; 14'h3E49: rddata <= 8'h00; 14'h3E4A: rddata <= 8'h3F; 14'h3E4B: rddata <= 8'h30;
            14'h3E4C: rddata <= 8'h37; 14'h3E4D: rddata <= 8'h36; 14'h3E4E: rddata <= 8'h36; 14'h3E4F: rddata <= 8'h36;
            14'h3E50: rddata <= 8'h36; 14'h3E51: rddata <= 8'h36; 14'h3E52: rddata <= 8'hF7; 14'h3E53: rddata <= 8'h00;
            14'h3E54: rddata <= 8'hFF; 14'h3E55: rddata <= 8'h00; 14'h3E56: rddata <= 8'h00; 14'h3E57: rddata <= 8'h00;
            14'h3E58: rddata <= 8'h00; 14'h3E59: rddata <= 8'h00; 14'h3E5A: rddata <= 8'hFF; 14'h3E5B: rddata <= 8'h00;
            14'h3E5C: rddata <= 8'hF7; 14'h3E5D: rddata <= 8'h36; 14'h3E5E: rddata <= 8'h36; 14'h3E5F: rddata <= 8'h36;
            14'h3E60: rddata <= 8'h36; 14'h3E61: rddata <= 8'h36; 14'h3E62: rddata <= 8'h37; 14'h3E63: rddata <= 8'h30;
            14'h3E64: rddata <= 8'h37; 14'h3E65: rddata <= 8'h36; 14'h3E66: rddata <= 8'h36; 14'h3E67: rddata <= 8'h36;
            14'h3E68: rddata <= 8'h00; 14'h3E69: rddata <= 8'h00; 14'h3E6A: rddata <= 8'hFF; 14'h3E6B: rddata <= 8'h00;
            14'h3E6C: rddata <= 8'hFF; 14'h3E6D: rddata <= 8'h00; 14'h3E6E: rddata <= 8'h00; 14'h3E6F: rddata <= 8'h00;
            14'h3E70: rddata <= 8'h36; 14'h3E71: rddata <= 8'h36; 14'h3E72: rddata <= 8'hF7; 14'h3E73: rddata <= 8'h00;
            14'h3E74: rddata <= 8'hF7; 14'h3E75: rddata <= 8'h36; 14'h3E76: rddata <= 8'h36; 14'h3E77: rddata <= 8'h36;
            14'h3E78: rddata <= 8'h18; 14'h3E79: rddata <= 8'h18; 14'h3E7A: rddata <= 8'hFF; 14'h3E7B: rddata <= 8'h00;
            14'h3E7C: rddata <= 8'hFF; 14'h3E7D: rddata <= 8'h00; 14'h3E7E: rddata <= 8'h00; 14'h3E7F: rddata <= 8'h00;
            14'h3E80: rddata <= 8'h36; 14'h3E81: rddata <= 8'h36; 14'h3E82: rddata <= 8'h36; 14'h3E83: rddata <= 8'h36;
            14'h3E84: rddata <= 8'hFF; 14'h3E85: rddata <= 8'h00; 14'h3E86: rddata <= 8'h00; 14'h3E87: rddata <= 8'h00;
            14'h3E88: rddata <= 8'h00; 14'h3E89: rddata <= 8'h00; 14'h3E8A: rddata <= 8'hFF; 14'h3E8B: rddata <= 8'h00;
            14'h3E8C: rddata <= 8'hFF; 14'h3E8D: rddata <= 8'h18; 14'h3E8E: rddata <= 8'h18; 14'h3E8F: rddata <= 8'h18;
            14'h3E90: rddata <= 8'h00; 14'h3E91: rddata <= 8'h00; 14'h3E92: rddata <= 8'h00; 14'h3E93: rddata <= 8'h00;
            14'h3E94: rddata <= 8'hFF; 14'h3E95: rddata <= 8'h36; 14'h3E96: rddata <= 8'h36; 14'h3E97: rddata <= 8'h36;
            14'h3E98: rddata <= 8'h36; 14'h3E99: rddata <= 8'h36; 14'h3E9A: rddata <= 8'h36; 14'h3E9B: rddata <= 8'h36;
            14'h3E9C: rddata <= 8'h3F; 14'h3E9D: rddata <= 8'h00; 14'h3E9E: rddata <= 8'h00; 14'h3E9F: rddata <= 8'h00;
            14'h3EA0: rddata <= 8'h18; 14'h3EA1: rddata <= 8'h18; 14'h3EA2: rddata <= 8'h1F; 14'h3EA3: rddata <= 8'h18;
            14'h3EA4: rddata <= 8'h1F; 14'h3EA5: rddata <= 8'h00; 14'h3EA6: rddata <= 8'h00; 14'h3EA7: rddata <= 8'h00;
            14'h3EA8: rddata <= 8'h00; 14'h3EA9: rddata <= 8'h00; 14'h3EAA: rddata <= 8'h1F; 14'h3EAB: rddata <= 8'h18;
            14'h3EAC: rddata <= 8'h1F; 14'h3EAD: rddata <= 8'h18; 14'h3EAE: rddata <= 8'h18; 14'h3EAF: rddata <= 8'h18;
            14'h3EB0: rddata <= 8'h00; 14'h3EB1: rddata <= 8'h00; 14'h3EB2: rddata <= 8'h00; 14'h3EB3: rddata <= 8'h00;
            14'h3EB4: rddata <= 8'h3F; 14'h3EB5: rddata <= 8'h36; 14'h3EB6: rddata <= 8'h36; 14'h3EB7: rddata <= 8'h36;
            14'h3EB8: rddata <= 8'h36; 14'h3EB9: rddata <= 8'h36; 14'h3EBA: rddata <= 8'h36; 14'h3EBB: rddata <= 8'h36;
            14'h3EBC: rddata <= 8'hFF; 14'h3EBD: rddata <= 8'h36; 14'h3EBE: rddata <= 8'h36; 14'h3EBF: rddata <= 8'h36;
            14'h3EC0: rddata <= 8'h18; 14'h3EC1: rddata <= 8'h18; 14'h3EC2: rddata <= 8'hFF; 14'h3EC3: rddata <= 8'h18;
            14'h3EC4: rddata <= 8'hFF; 14'h3EC5: rddata <= 8'h18; 14'h3EC6: rddata <= 8'h18; 14'h3EC7: rddata <= 8'h18;
            14'h3EC8: rddata <= 8'h18; 14'h3EC9: rddata <= 8'h18; 14'h3ECA: rddata <= 8'h18; 14'h3ECB: rddata <= 8'h18;
            14'h3ECC: rddata <= 8'hF8; 14'h3ECD: rddata <= 8'h00; 14'h3ECE: rddata <= 8'h00; 14'h3ECF: rddata <= 8'h00;
            14'h3ED0: rddata <= 8'h00; 14'h3ED1: rddata <= 8'h00; 14'h3ED2: rddata <= 8'h00; 14'h3ED3: rddata <= 8'h00;
            14'h3ED4: rddata <= 8'h1F; 14'h3ED5: rddata <= 8'h18; 14'h3ED6: rddata <= 8'h18; 14'h3ED7: rddata <= 8'h18;
            14'h3ED8: rddata <= 8'hFF; 14'h3ED9: rddata <= 8'hFF; 14'h3EDA: rddata <= 8'hFF; 14'h3EDB: rddata <= 8'hFF;
            14'h3EDC: rddata <= 8'hFF; 14'h3EDD: rddata <= 8'hFF; 14'h3EDE: rddata <= 8'hFF; 14'h3EDF: rddata <= 8'hFF;
            14'h3EE0: rddata <= 8'h00; 14'h3EE1: rddata <= 8'h00; 14'h3EE2: rddata <= 8'h00; 14'h3EE3: rddata <= 8'h00;
            14'h3EE4: rddata <= 8'hFF; 14'h3EE5: rddata <= 8'hFF; 14'h3EE6: rddata <= 8'hFF; 14'h3EE7: rddata <= 8'hFF;
            14'h3EE8: rddata <= 8'hF0; 14'h3EE9: rddata <= 8'hF0; 14'h3EEA: rddata <= 8'hF0; 14'h3EEB: rddata <= 8'hF0;
            14'h3EEC: rddata <= 8'hF0; 14'h3EED: rddata <= 8'hF0; 14'h3EEE: rddata <= 8'hF0; 14'h3EEF: rddata <= 8'hF0;
            14'h3EF0: rddata <= 8'h0F; 14'h3EF1: rddata <= 8'h0F; 14'h3EF2: rddata <= 8'h0F; 14'h3EF3: rddata <= 8'h0F;
            14'h3EF4: rddata <= 8'h0F; 14'h3EF5: rddata <= 8'h0F; 14'h3EF6: rddata <= 8'h0F; 14'h3EF7: rddata <= 8'h0F;
            14'h3EF8: rddata <= 8'hFF; 14'h3EF9: rddata <= 8'hFF; 14'h3EFA: rddata <= 8'hFF; 14'h3EFB: rddata <= 8'hFF;
            14'h3EFC: rddata <= 8'h00; 14'h3EFD: rddata <= 8'h00; 14'h3EFE: rddata <= 8'h00; 14'h3EFF: rddata <= 8'h00;
            14'h3F00: rddata <= 8'h00; 14'h3F01: rddata <= 8'h00; 14'h3F02: rddata <= 8'h3B; 14'h3F03: rddata <= 8'h6E;
            14'h3F04: rddata <= 8'h64; 14'h3F05: rddata <= 8'h6E; 14'h3F06: rddata <= 8'h3B; 14'h3F07: rddata <= 8'h00;
            14'h3F08: rddata <= 8'h3C; 14'h3F09: rddata <= 8'h66; 14'h3F0A: rddata <= 8'h66; 14'h3F0B: rddata <= 8'h6C;
            14'h3F0C: rddata <= 8'h63; 14'h3F0D: rddata <= 8'h63; 14'h3F0E: rddata <= 8'h66; 14'h3F0F: rddata <= 8'h00;
            14'h3F10: rddata <= 8'h7E; 14'h3F11: rddata <= 8'h66; 14'h3F12: rddata <= 8'h60; 14'h3F13: rddata <= 8'h60;
            14'h3F14: rddata <= 8'h60; 14'h3F15: rddata <= 8'h60; 14'h3F16: rddata <= 8'h60; 14'h3F17: rddata <= 8'h00;
            14'h3F18: rddata <= 8'h00; 14'h3F19: rddata <= 8'h7F; 14'h3F1A: rddata <= 8'h36; 14'h3F1B: rddata <= 8'h36;
            14'h3F1C: rddata <= 8'h36; 14'h3F1D: rddata <= 8'h36; 14'h3F1E: rddata <= 8'h36; 14'h3F1F: rddata <= 8'h00;
            14'h3F20: rddata <= 8'h7E; 14'h3F21: rddata <= 8'h66; 14'h3F22: rddata <= 8'h30; 14'h3F23: rddata <= 8'h18;
            14'h3F24: rddata <= 8'h30; 14'h3F25: rddata <= 8'h66; 14'h3F26: rddata <= 8'h7E; 14'h3F27: rddata <= 8'h00;
            14'h3F28: rddata <= 8'h00; 14'h3F29: rddata <= 8'h00; 14'h3F2A: rddata <= 8'h3F; 14'h3F2B: rddata <= 8'h6C;
            14'h3F2C: rddata <= 8'h6C; 14'h3F2D: rddata <= 8'h6C; 14'h3F2E: rddata <= 8'h38; 14'h3F2F: rddata <= 8'h00;
            14'h3F30: rddata <= 8'h00; 14'h3F31: rddata <= 8'h33; 14'h3F32: rddata <= 8'h33; 14'h3F33: rddata <= 8'h33;
            14'h3F34: rddata <= 8'h33; 14'h3F35: rddata <= 8'h3E; 14'h3F36: rddata <= 8'h30; 14'h3F37: rddata <= 8'h60;
            14'h3F38: rddata <= 8'h00; 14'h3F39: rddata <= 8'h3B; 14'h3F3A: rddata <= 8'h6E; 14'h3F3B: rddata <= 8'h0C;
            14'h3F3C: rddata <= 8'h0C; 14'h3F3D: rddata <= 8'h0C; 14'h3F3E: rddata <= 8'h0C; 14'h3F3F: rddata <= 8'h00;
            14'h3F40: rddata <= 8'h7E; 14'h3F41: rddata <= 8'h18; 14'h3F42: rddata <= 8'h3C; 14'h3F43: rddata <= 8'h66;
            14'h3F44: rddata <= 8'h66; 14'h3F45: rddata <= 8'h3C; 14'h3F46: rddata <= 8'h18; 14'h3F47: rddata <= 8'h7E;
            14'h3F48: rddata <= 8'h1C; 14'h3F49: rddata <= 8'h36; 14'h3F4A: rddata <= 8'h63; 14'h3F4B: rddata <= 8'h7F;
            14'h3F4C: rddata <= 8'h63; 14'h3F4D: rddata <= 8'h36; 14'h3F4E: rddata <= 8'h1C; 14'h3F4F: rddata <= 8'h00;
            14'h3F50: rddata <= 8'h1C; 14'h3F51: rddata <= 8'h36; 14'h3F52: rddata <= 8'h63; 14'h3F53: rddata <= 8'h63;
            14'h3F54: rddata <= 8'h36; 14'h3F55: rddata <= 8'h36; 14'h3F56: rddata <= 8'h77; 14'h3F57: rddata <= 8'h00;
            14'h3F58: rddata <= 8'h0E; 14'h3F59: rddata <= 8'h18; 14'h3F5A: rddata <= 8'h0C; 14'h3F5B: rddata <= 8'h3E;
            14'h3F5C: rddata <= 8'h66; 14'h3F5D: rddata <= 8'h66; 14'h3F5E: rddata <= 8'h3C; 14'h3F5F: rddata <= 8'h00;
            14'h3F60: rddata <= 8'h00; 14'h3F61: rddata <= 8'h00; 14'h3F62: rddata <= 8'h7E; 14'h3F63: rddata <= 8'hDB;
            14'h3F64: rddata <= 8'hDB; 14'h3F65: rddata <= 8'h7E; 14'h3F66: rddata <= 8'h00; 14'h3F67: rddata <= 8'h00;
            14'h3F68: rddata <= 8'h06; 14'h3F69: rddata <= 8'h0C; 14'h3F6A: rddata <= 8'h7E; 14'h3F6B: rddata <= 8'hDB;
            14'h3F6C: rddata <= 8'hDB; 14'h3F6D: rddata <= 8'h7E; 14'h3F6E: rddata <= 8'h60; 14'h3F6F: rddata <= 8'hC0;
            14'h3F70: rddata <= 8'h1C; 14'h3F71: rddata <= 8'h30; 14'h3F72: rddata <= 8'h60; 14'h3F73: rddata <= 8'h7C;
            14'h3F74: rddata <= 8'h60; 14'h3F75: rddata <= 8'h30; 14'h3F76: rddata <= 8'h1C; 14'h3F77: rddata <= 8'h00;
            14'h3F78: rddata <= 8'h3C; 14'h3F79: rddata <= 8'h66; 14'h3F7A: rddata <= 8'h66; 14'h3F7B: rddata <= 8'h66;
            14'h3F7C: rddata <= 8'h66; 14'h3F7D: rddata <= 8'h66; 14'h3F7E: rddata <= 8'h66; 14'h3F7F: rddata <= 8'h00;
            14'h3F80: rddata <= 8'h00; 14'h3F81: rddata <= 8'h7E; 14'h3F82: rddata <= 8'h00; 14'h3F83: rddata <= 8'h7E;
            14'h3F84: rddata <= 8'h00; 14'h3F85: rddata <= 8'h7E; 14'h3F86: rddata <= 8'h00; 14'h3F87: rddata <= 8'h00;
            14'h3F88: rddata <= 8'h18; 14'h3F89: rddata <= 8'h18; 14'h3F8A: rddata <= 8'h7E; 14'h3F8B: rddata <= 8'h18;
            14'h3F8C: rddata <= 8'h18; 14'h3F8D: rddata <= 8'h00; 14'h3F8E: rddata <= 8'h7E; 14'h3F8F: rddata <= 8'h00;
            14'h3F90: rddata <= 8'h30; 14'h3F91: rddata <= 8'h18; 14'h3F92: rddata <= 8'h0C; 14'h3F93: rddata <= 8'h18;
            14'h3F94: rddata <= 8'h30; 14'h3F95: rddata <= 8'h00; 14'h3F96: rddata <= 8'h7E; 14'h3F97: rddata <= 8'h00;
            14'h3F98: rddata <= 8'h0C; 14'h3F99: rddata <= 8'h18; 14'h3F9A: rddata <= 8'h30; 14'h3F9B: rddata <= 8'h18;
            14'h3F9C: rddata <= 8'h0C; 14'h3F9D: rddata <= 8'h00; 14'h3F9E: rddata <= 8'h7E; 14'h3F9F: rddata <= 8'h00;
            14'h3FA0: rddata <= 8'h0E; 14'h3FA1: rddata <= 8'h1B; 14'h3FA2: rddata <= 8'h1B; 14'h3FA3: rddata <= 8'h18;
            14'h3FA4: rddata <= 8'h18; 14'h3FA5: rddata <= 8'h18; 14'h3FA6: rddata <= 8'h18; 14'h3FA7: rddata <= 8'h18;
            14'h3FA8: rddata <= 8'h18; 14'h3FA9: rddata <= 8'h18; 14'h3FAA: rddata <= 8'h18; 14'h3FAB: rddata <= 8'h18;
            14'h3FAC: rddata <= 8'h18; 14'h3FAD: rddata <= 8'hD8; 14'h3FAE: rddata <= 8'hD8; 14'h3FAF: rddata <= 8'h70;
            14'h3FB0: rddata <= 8'h18; 14'h3FB1: rddata <= 8'h18; 14'h3FB2: rddata <= 8'h00; 14'h3FB3: rddata <= 8'h7E;
            14'h3FB4: rddata <= 8'h00; 14'h3FB5: rddata <= 8'h18; 14'h3FB6: rddata <= 8'h18; 14'h3FB7: rddata <= 8'h00;
            14'h3FB8: rddata <= 8'h00; 14'h3FB9: rddata <= 8'h76; 14'h3FBA: rddata <= 8'hDC; 14'h3FBB: rddata <= 8'h00;
            14'h3FBC: rddata <= 8'h76; 14'h3FBD: rddata <= 8'hDC; 14'h3FBE: rddata <= 8'h00; 14'h3FBF: rddata <= 8'h00;
            14'h3FC0: rddata <= 8'h38; 14'h3FC1: rddata <= 8'h6C; 14'h3FC2: rddata <= 8'h6C; 14'h3FC3: rddata <= 8'h38;
            14'h3FC4: rddata <= 8'h00; 14'h3FC5: rddata <= 8'h00; 14'h3FC6: rddata <= 8'h00; 14'h3FC7: rddata <= 8'h00;
            14'h3FC8: rddata <= 8'h00; 14'h3FC9: rddata <= 8'h00; 14'h3FCA: rddata <= 8'h00; 14'h3FCB: rddata <= 8'h18;
            14'h3FCC: rddata <= 8'h18; 14'h3FCD: rddata <= 8'h00; 14'h3FCE: rddata <= 8'h00; 14'h3FCF: rddata <= 8'h00;
            14'h3FD0: rddata <= 8'h00; 14'h3FD1: rddata <= 8'h00; 14'h3FD2: rddata <= 8'h00; 14'h3FD3: rddata <= 8'h00;
            14'h3FD4: rddata <= 8'h18; 14'h3FD5: rddata <= 8'h00; 14'h3FD6: rddata <= 8'h00; 14'h3FD7: rddata <= 8'h00;
            14'h3FD8: rddata <= 8'h0F; 14'h3FD9: rddata <= 8'h0C; 14'h3FDA: rddata <= 8'h0C; 14'h3FDB: rddata <= 8'h0C;
            14'h3FDC: rddata <= 8'hEC; 14'h3FDD: rddata <= 8'h6C; 14'h3FDE: rddata <= 8'h3C; 14'h3FDF: rddata <= 8'h1C;
            14'h3FE0: rddata <= 8'h78; 14'h3FE1: rddata <= 8'h6C; 14'h3FE2: rddata <= 8'h6C; 14'h3FE3: rddata <= 8'h6C;
            14'h3FE4: rddata <= 8'h6C; 14'h3FE5: rddata <= 8'h00; 14'h3FE6: rddata <= 8'h00; 14'h3FE7: rddata <= 8'h00;
            14'h3FE8: rddata <= 8'h38; 14'h3FE9: rddata <= 8'h0C; 14'h3FEA: rddata <= 8'h18; 14'h3FEB: rddata <= 8'h30;
            14'h3FEC: rddata <= 8'h3C; 14'h3FED: rddata <= 8'h00; 14'h3FEE: rddata <= 8'h00; 14'h3FEF: rddata <= 8'h00;
            14'h3FF0: rddata <= 8'h00; 14'h3FF1: rddata <= 8'h00; 14'h3FF2: rddata <= 8'h3C; 14'h3FF3: rddata <= 8'h3C;
            14'h3FF4: rddata <= 8'h3C; 14'h3FF5: rddata <= 8'h3C; 14'h3FF6: rddata <= 8'h00; 14'h3FF7: rddata <= 8'h00;
            14'h3FF8: rddata <= 8'h00; 14'h3FF9: rddata <= 8'h00; 14'h3FFA: rddata <= 8'h00; 14'h3FFB: rddata <= 8'h00;
            14'h3FFC: rddata <= 8'h00; 14'h3FFD: rddata <= 8'h00; 14'h3FFE: rddata <= 8'h00; 14'h3FFF: rddata <= 8'h00;
        endcase

endmodule
