module videoram(
    // First port - CPU access
    input  wire        p1_clk,
    input  wire [10:0] p1_addr,
    output wire  [7:0] p1_rddata,
    input  wire  [7:0] p1_wrdata,
    input  wire        p1_wren,

    // Second port - Video access
    input  wire        p2_clk,
    input  wire  [9:0] p2_addr,
    output wire [15:0] p2_rddata);

    RAMB16_S9_S18 #(
        .INIT_A(9'h000),                // Value of output RAM registers on Port A at startup
        .INIT_B(18'h00000),             // Value of output RAM registers on Port B at startup
        .SRVAL_A(9'h000),               // Port A output value upon SSR assertion
        .SRVAL_B(18'h00000),            // Port B output value upon SSR assertion
        .WRITE_MODE_A("WRITE_FIRST"),   // WRITE_FIRST, READ_FIRST or NO_CHANGE
        .WRITE_MODE_B("WRITE_FIRST"),   // WRITE_FIRST, READ_FIRST or NO_CHANGE
        .SIM_COLLISION_CHECK("NONE"),   // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL"

        // The following INIT_xx declarations specify the initial contents of the RAM
        // Port A Address 0 to 511, Port B Address 0 to 255
        .INIT_00(256'hE420E420E420E420E420E420E420E420E420E420E420E420E420E420E420DED8),
        .INIT_01(256'hE420E420E420E420E420E420E420E420E420E420E420E420E420E420E420E420),
        .INIT_02(256'hE420E420E420E420E420E420E420E420E420E420E420E420E420E420E420E420),
        .INIT_03(256'hE420E42074C6E420E420E420E420E420E420E420E420E420E420E420E420E420),
        .INIT_04(256'hE420E42074C6E420E420E420E420E420E420E420E42074D174D084D174D0E420),
        .INIT_05(256'hE420E420E42074C4E420E420E420E42074C6E420E420E420E420E42074C6E420),
        .INIT_06(256'h74C6E420E420EED2EED2E0910E81E420E420E420E420E420E42074C6E420E420),
        .INIT_07(256'hE420E420E42034D234D2E420E420E42074C6E420E420E420E420E420E420E420),
        .INIT_08(256'h04DD04DC048D0418048D0418048D0418048D0418E420E420E420E420E420E420),
        .INIT_09(256'hE420E420E420E420E420E420E420E420E420E420E420EED2EED2E0910E81E420),
        .INIT_0A(256'h87D087D087D074C0E420E420E420E420E420E42034DBC47FC47F34CBE420E420),
        .INIT_0B(256'h87D087D087D07EC0EED2E0910E8187D087D087D087D087D087D087D087D087D0),
        .INIT_0C(256'h74C6E42034DBC47FC47F34CBE420E420E420E420E42074C6E420E420E4C1E7C0),
        .INIT_0D(256'h7F7F7F7F872E7F7F7F7F7F7F7F7F7F7F87C67F7F87D087D074C0E420E420E420),
        .INIT_0E(256'hE420E420E420E420E420E4C1EF7FEF7FE7C07F7F7F7F7F7F7EC0E0910E817F7F),
        .INIT_0F(256'h7F7F7F7F7F7F87D087D074C0E420E420E420E420E42034C234C2E420E420E420),

        // Port A Address 512 to 1023, Port B Address 256 to 511
        .INIT_10(256'hEF7FE7C07F7F7F7F872E7F7F7F7F7F7F87C67F7F7F7F7F7F7F7F872E7F7F87C6),
        .INIT_11(256'hE420E420E420E420E420E420E420E42074C6E42074C4E420E4C1EF7FF01FF01F),
        .INIT_12(256'h7F7F872E7F7F7F7F87C67F7F7F7F7F7F7F7F872E7F7F7F7F87D087D074C0E420),
        .INIT_13(256'hE420E420E420E4C1EF7FEF7F0F1F0F1FEF7FEF7FE7C07F7F7F7F7F7F872E7F7F),
        .INIT_14(256'h7F7F872E872E7F7F7F7F87D087D074C0E420E420E42074C4E420E420E420E420),
        .INIT_15(256'hEF7FEF7FEF7FE7C07F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F),
        .INIT_16(256'hE420E420E420E420E420E420E420E420E420E420E4C1EF7FEF7FEF7FEF7FEF7F),
        .INIT_17(256'hE080E080E080E7C07F7FE7C1E0807EC2E080E0807EC27EC2E080E080E0800E97),
        .INIT_18(256'hE420E420EB917E6B7E437E697E4EEF7F7E747E53EF7F0E97E0807EC27EC27EC2),
        .INIT_19(256'h0E900E900E90EF7FEF7FEF7FEF7F0E97E420E420E420E42014D4E420E42074C6),
        .INIT_1A(256'h0E90EF7FEF7F0E97EF7FEF7F0E900E900E90EF7FEF7FEF7F7EC2EF7FEF7FEF7F),
        .INIT_1B(256'hE420E420E420E42034C8E420E420E42074C4E420E091EF7F0E900E900E900E90),
        .INIT_1C(256'hC7D1E091EF7FEF7F1E5EEF7FEF7F0E81C7D1C7D1C7D1E091EF7FEF7FEF7F0E97),
        .INIT_1D(256'hE420E420E0910E810CC97CD00C8F7CD00CD7E091EF7F0E97EF7F0E81C7D1C7D1),
        .INIT_1E(256'h7CD07CD07CD0E091EF7FEF7FEF7F0E97E420E420E42024C112C624C0E420E420),
        .INIT_1F(256'h7CD0E091EF7F0E97EF7F0E817CD07CD07CD0E091EF7F1E7BDED31E7DEF7F0E81),

        // Port A Address 1024 to 1535, Port B Address 512 to 767
        .INIT_20(256'hE420E42024C142C6227F12C424C0E420E420E420E0910E817CD00C9D0C080C9C),
        .INIT_21(256'h1C96E091EF7FE0AFE0AFE0AFEF7F0E81DC195CDC5C9EE091EF7FEF7FEF7F0E97),
        .INIT_22(256'hE42074C6E0910E817CD00CC90C120CD77CD0E091EF7F0E97EF7F0E817CD04C0E),
        .INIT_23(256'hE080E080E080EF7FEF7FEF7FEF7F0E9774C6E42024C1247F12C672C624C0E420),
        .INIT_24(256'hE080EF7FEF7F0E97EF7FEF7FE080E080E080EF7F0E99C7D17CD7C7D1E099EF7F),
        .INIT_25(256'hE420E42024C152C4227F227F24C0E420E42064C96E896ED7E080E080E080E080),
        .INIT_26(256'hEF7FEF7F0E997CD01C8F7CD0E099EF7FEF7FEF7FEF7FEF7FEF7FEF7FEF7F0E97),
        .INIT_27(256'hE420E4207E96EF7FEF7FEF7FEF7FEF7FEF7F7ED27ED20E97EF7FEF7FEF7FEF7F),
        .INIT_28(256'hEF7FEF7FEF7F7ED27E20EF7FEF7F0E97E420E42024C1247F32C642C624C0E420),
        .INIT_29(256'h7EC10720072007207EC0EF7FEF7FEF7FEF7FEF7F0E997CD01C927CD0E099EF7F),
        .INIT_2A(256'h74D2E420E420E420E486E420E42074C1E4C674DBD7C27ECBEF7FEF7FEF7FEF7F),
        .INIT_2B(256'hEF7FEF7F0E997CD0FC147CD0E099EF7F7EC57ED27EC1072007207EC07ED20E97),
        .INIT_2C(256'hE42074C107207EC0EF7FEF7F7ED27EC107200720872E072007207EC0EF7F7ED2),
        .INIT_2D(256'h072007200720072087C6072007200720072007200720072087C60720072087C6),
        .INIT_2E(256'h07200720072007200720072007200720072078C08F7F8F7F8F7F08208F7F87C0),
        .INIT_2F(256'h072087C6072007200720872E87C6072007200720072007200720072007200720),

        // Port A Address 1536 to 2047, Port B Address 768 to 1023
        .INIT_30(256'h87C6072078C08F7F8F7F082008208F7F87C0072087C6072007208720872E0720),
        .INIT_31(256'h87C60720072087C60720872E072087C60720072087C60720872E072087C60720),
        .INIT_32(256'h082087C00720872E072007200720072087C6072087C60720072087C607200720),
        .INIT_33(256'h0720872E07200720072087C60720072007200720072078C08F7F082008200820),
        .INIT_34(256'h072087C607200720072007200720872E072007200720072087C607200720872E),
        .INIT_35(256'h87C60720872E072078C08F7F0820082008208F7F87C00720072087C607200720),
        .INIT_36(256'h0720872E07200720072007200720072087C60720072007200720072007200720),
        .INIT_37(256'h0820082058EC8F898F898F898F898F898F898F898F898F898F898F898F898F89),
        .INIT_38(256'h8F898F898F898F898F898F898F898F898F898F898F898F898F898F7F28150820),
        .INIT_39(256'h0820082038AC0820082038AC082048198F898F898F898F898F898F898F898F89),
        .INIT_3A(256'h38AC0820082038AC08200820D8180820082038AC0820082038AC0820082038AC),
        .INIT_3B(256'h082038AC0820082038AC0820082038AC0820082038AC0820D89A38AC08200820),
        .INIT_3C(256'h08200820082008200820082008200820D89B0820082008200820082008200820),
        .INIT_3D(256'h0820082008200820082008200820082008200820188708200820082008200820),
        .INIT_3E(256'h0000000000000000000000000000000008200820082048190820082008200820),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),

        // The next set of INITP_xx are for the parity bits
        // Port A Address 0 to 511, Port B Address 0 to 255
        .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        // Port A Address 512 to 1023, Port B Address 256 to 511
        .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        // Port A Address 1024 to 1535, Port B Address 512 to 767
        .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        // Port A Address 1536 to 2047, Port B Address 768 to 1024
        .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000))
    
    RAMB16_S9_S18_inst(
        // Port-A
        .CLKA(p1_clk),      // Clock
        .SSRA(1'b0),        // Synchronous Set/Reset Input
        .ADDRA(p1_addr),    // 11-bit Address Input
        .DOA(p1_rddata),    // 8-bit Data Output
        .DOPA(),            // 1-bit Parity Output
        .DIA(p1_wrdata),    // 8-bit Data Input
        .DIPA(1'b0),        // 1-bit parity Input
        .ENA(1'b1),         // RAM Enable Input
        .WEA(p1_wren),      // Write Enable Input

        // Port-B
        .CLKB(p2_clk),      // Clock
        .SSRB(1'b0),        // Synchronous Set/Reset Input
        .ADDRB(p2_addr),    // 10-bit Address Input
        .DOB(p2_rddata),    // 16-bit Data Output
        .DOPB(),            // 2-bit Parity Output
        .DIB(16'b0),        // 16-bit Data Input
        .DIPB(2'b0),        // 2-bit parity Input
        .ENB(1'b1),         // RAM Enable Input
        .WEB(1'b0)          // Write Enable Input
    );

endmodule
