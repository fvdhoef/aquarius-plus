module rom(
    input  wire        clk,
    input  wire [15:0] addr,
    output reg   [7:0] rddata);

    reg addr_r;
    always @(posedge clk) addr_r <= addr;

    wire [7:0] rddata_00;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000198AC30670C3D03AFE7E2303C4C2E323BEE37E000B2206822000C3),
        .INIT_01(256'hD9E523E1D93803C30000E9DD38062ADDC914EBC2B738E73A0000C9937DC0927C),
        .INIT_02(256'h21E01111385D222FFF21FFD3AF1D94CD073E203638012A1D94CD0B3E38A031C9),
        .INIT_03(256'hC3380932FFD3AEFA20058023860C06EB1920B77EF628BE830F0F1A231B1B0081),
        .INIT_04(256'h06B0ED00190100B521321011B0ED00050100B02131A111002C332424372B2006),
        .INIT_05(256'h52555445522073736572504349534142EF1800CFCD060600CFCD020600CFCD03),
        .INIT_06(256'hFE1E80CD400021F92038FE7C2370340021007472617473206F742079656B204E),
        .INIT_07(256'h0187211A40CD0BE5CDFFD338093A1D72CD0B3EC9F020B57C2B062803FE1A280D),
        .INIT_08(256'h712F7E772F4677A90B28B57C4E232003C339003238A932AFB0ED380311005101),
        .INIT_09(256'hE5CD3865311FF2CD0BBECD384B221938AD22FFCE110BB7DAE73A2C112BEF28B8),
        .INIT_0A(256'h0B0402C3380932FFD3AF175FEDF418132B0420BE1FE8CAB71A0082112005210B),
        .INIT_0B(256'h6E492074666F736F7263694D2079622032383931200520746867697279706F43),
        .INIT_0C(256'h3E4700DE786700DE7C6F00D6000020000000A300003B0697C3000A3253202E63),
        .INIT_0D(256'hCDBC65989F1A0A9999D1539847DD0A98B3952298761C3999CA4A35000000C900),
        .INIT_0E(256'hCC0893071C0D1305BC0C213901FFFE3964000E28000000804FC752983E77D698),
        .INIT_0F(256'hBC0B6D0B3B1B1507B507800C1F071E06F806CB0C05079C06BE06DC073108BE10),
        .INIT_10(256'h2E10A83803150915B114F50BBD1AD61A4C1A4F1C081C2C0CCD0567056C0C4B07),
        .INIT_11(256'h211013100210840E290FF30B631985197018DD18D717CD1385186617750B330B),
        .INIT_12(256'hCC444145D24D49C45455504EC9415441C4545845CE524FC6444EC51059105010),
        .INIT_13(256'h4D45D24E52555445D24255534FC745524F545345D246C94E55D24F544FC75445),
        .INIT_14(256'h544E4FC3544E4952D0454B4FD04645C459504FC3544E495250CC4ECF504F54D3),
        .INIT_15(256'h534552D0544553D045564153C344414F4CC35241454CC35453494CCC545349CC),
        .INIT_16(256'h4E4548D42459454B4EC9284350D34EC64FD4284241D45745CE444E554FD35445),
        .INIT_17(256'h5253D55342C1544EC94E47D3BCBDBE52CF444EC1DEAFAAADAB504554D3544FCE),
        .INIT_18(256'hC14E41D44E49D3534FC35058C5474FCC444ED25251D3534FD0534F50CC4552C6),
        .INIT_19(256'h484749D224544645CC245248C34353C14C41D6245254D34E45CC4B4545D04E54),
        .INIT_1A(256'hA8460AA950177E7F142D7C13C97C125C79165C7980544E494FD0244449CD2454),
        .INIT_1B(256'h4F47524E53464E006B61657242000A0D6B4F00206E69200007726F727245200A),
        .INIT_1C(256'h214F4D46554E435453534C534F4D544449302F444453424C554D4F564F434644),
        .INIT_1D(256'hC92AE51809C8E1000D01E7EB0228EBB37A6960E52346234EC081FE237E390004),
        .INIT_1E(256'h00F70BE5CD181E01241E010A1E01221E01121E01001E01141E01021E384D2238),
        .INIT_1F(256'h166DC43CA57C384D2A0E9DCD036121DFD7DF7EDF3F3E195701F703792119DECD),
        .INIT_20(256'hD7F5380D85CD384D22FFFF210E9DCD036E2119DECD380832AF19BECD02F7C13E),
        .INIT_21(256'h049FCDF5B7D738CC32AFC5D5064BD203F7F1D14704BCCDD5069CCDF5F0283D3C),
        .INIT_22(256'h2A2128F1D138D6226960F920E71303021A38D62AEB1030C5B706F3CAF5F10638),
        .INIT_23(256'hF920B71323771A386011237223732323D174EB38D622E10B92CDE509C1E338D6),
        .INIT_24(256'h2AEA18722373EBFC2023BEAF2323230414CAB6237E6B62EB2305F70BCBCD04F7),
        .INIT_25(256'h38AC32AFE618D03FC83F6F66237E6960E76F66237E2323C82BB6237E4D44384F),
        .INIT_26(256'h3E3FFE053CC27EB738AC3A055ECAB70558CA22FE47053CCA20FE7E386011050E),
        .INIT_27(256'h7BFE073861FE7E7F06C5053601C5024411D5053CDA3CFE053830FE7E053CCA95),
        .INIT_28(256'h88FE784F0532FAB71A13E5EBF320B9C87FE67E040507F2B623EB4E775FE60330),
        .INIT_29(256'h0C131223D1C179EB0AF7C9EBF148D318E1E728B95FE6023861FE7E232BD70220),
        .INIT_2A(256'h5F21F318130C1223E428B80928B77E4704C5C254D638AC32032049FE04283AD6),
        .INIT_2B(256'h782346234EE1C5049FCDC1C0069CCD380832173E384732013EC9121312131238),
        .INIT_2C(256'h0597F2DD28B7237EDFE1203E1675CDEBE52356235E19EACDC51A25CD0402CAB1),
        .INIT_2D(256'hCB32643EDC1805B1F2B7131ADF7FE6F7200D05A8F2B7131A0245114F7FD616F7),
        .INIT_2E(256'hC72AE523235E2B562BD509142003A3CD3900022138C722071CCDE5C10731CD38),
        .INIT_2F(256'hCDA1CF0975CDE3384D2AE5E338C72AE50BA0CD080EEBD10CF9D1EA20D1E1E738),
        .INIT_30(256'hC5E1EF152ECDE50972CDD70A20013EA7FE7E5A51810001D5C5E1152ECDE50972),
        .INIT_31(256'hCAB6237E2303C4C2B714283AFE7E1FC2CD38CE2233C58106E338CE2AE533F5D5),
        .INIT_32(256'h064F0703C4D217F720FE0731DA80D6C8D5062C11D7EB384D22EB56235E230C29),
        .INIT_33(256'hFAEF0972CDD7C93D3C3F30FEF72820FED03AFE7E23EBC546234E0901D521EB00),
        .INIT_34(256'h0000112B03DBC3081EC851E1155BCDE50000119080011586DA90FE38E73A0697),
        .INIT_35(256'h18F7C9E1F1E518E1EB1900165F30D6F1291929196B621138E7199821F5E5D0D7),
        .INIT_36(256'hCD069CCDC533F58C3EE3384D2AE5E5C10BA0CD030E1018062C010BCFCD0BCBCA),
        .INIT_37(256'hFEF9039FCDFF16C003DBC30E1ED82B6960049FD404A2DCE1E7384D2AE523071E),
        .INIT_38(256'h000E3A01E13EE3062C210401C2B738CC3A0720B57C23384D22E103DBC2041E8C),
        .INIT_39(256'hE3F10985CDF538AB3AD5B0CF10D1CDF418F32822FE23C8B8C8B77E4748790006),
        .INIT_3A(256'h30D1E738DA2A0E30E7384F2A56235E2323E538E42AE50779CA0977CD1F38CE22),
        .INIT_3B(256'hC9E1D1153ACDE5C9E1153DCDE10FE4CD0E39CDEB0FE4CDD13E0930E738BD210F),
        .INIT_3C(256'h7E0985CDF318C02CFE069DCD0651CA780D4B2B88CF03288CFE477E0B54CD19F7),
        .INIT_3D(256'hEACC06F7D72B384732013E0650C306DCDAD7071ECAEF0975CD2BA5CF032888FE),
        .INIT_3E(256'h38AB3AE50985CDC10861CA3BFE44282CFEE5083ACAA3FE083ACAA0FE0866CA19),
        .INIT_3F(256'h38483A0D1884FE8638463A0828B738473A38E42A20360E5FCD1680CD0811C2B7)
    ) ram_00(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_00), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_01;
    RAMB16_S9_S9 #(
        .INIT_00(256'h38463A0828B738473AA318E10EA0C4AF0EA0CD19EAD4B83D8638003A09283C47),
        .INIT_01(256'h29CF0B53CDF520182FFC300ED60861D219EAD4B838003A4738493A082DC370FE),
        .INIT_02(256'h10DF203E473C0730832F38003A031838463A0853CAB738473A0F28E5A3D6F12B),
        .INIT_03(256'h000A0D7472617473206D6F7266206F6465523FC9384732AF07F707C1C3D7E1FD),
        .INIT_04(256'h08AAC2003E22FE7E0B45CD1AF70C01C30E9DCD086D21C103BEC2B738CD3A08F7),
        .INIT_05(256'h2AE505182C36071BCAC52BB77E230C26DAC10D5BCDE53E0EA0CDE53BCF0E60CD),
        .INIT_06(256'hCDDF3F3E0953C2B738CD3A1B282CFE7ED5E310D1CD2CCF01E338CD32AFF638DC),
        .INIT_07(256'h3A0C2822FE4757D71F28B738AB3A1CF7D5071BCAC5B72B7E230C26DAC1D10D5B),
        .INIT_08(256'hE1153ACDE315E5CDD7074AC3D5E3092021EB0E63CD2B2C063A16022857B738CD),
        .INIT_09(256'h0E9DC4094221B6D50C1AC2EBB738CD3AD108C9C2D72BE30880C22CFE0528D72B),
        .INIT_0A(256'hCA061EB6237E231120B7071CCD000A0D6465726F6E67692061727478453FC9E1),
        .INIT_0B(256'h03D9C3E8B78F38AB3A37F60985CD08F0C3E42083FED738C953ED56235E2303DB),
        .INIT_0C(256'h227E0975D478FE78C138D02A38D02209FDCD0BA0CD010ED500162B28CF01B0CF),
        .INIT_0D(256'h034C215F83070F7CCA7B3D38AB3A08205FA8D609E2D2AFFED0B2FED8A8FE38C3),
        .INIT_0E(256'hC338C32AC52346234E51581513CD4A43C5099401C50975CD23D0BA5678190016),
        .INIT_0F(256'hAF09F7E718D738C32203C4DA57BAAA1701FE0AD0D203FE0AD0DAAFD600160988),
        .INIT_10(256'h22FE0A3DCAA9FE15E5CA2EFEE928A8FE0A4ED20CC6CD15E5DA03D6CAD738AB32),
        .INIT_11(256'hCD7D16C929CF0983CD0A5FD2B2D60B40CAA2FE19FBCAA4FE0B05CAA6FE0E60CA),
        .INIT_12(256'hF7C9E11520CCB738AB3A38E422EBE510D1CDC9E10975CD150BCDE538D02A0988),
        .INIT_13(256'hEBE5E338E42AEB0976CD2CCF0983CD163829FE79D7C54F0700061A68CA18FE1B),
        .INIT_14(256'h14C82DFEC8A9FE15E96966234E09021501D50A4911E30A37CD0818E3EB0B54CD),
        .INIT_15(256'h79C1F10682CDF51523CDEBE3C1EBF10682CD0975CDF5AFF6C92BC8A8FEC82BFE),
        .INIT_16(256'hC3D0BA7864165F177A1F38AB3A0AE221E9B2784FB3E9A2784FA30ACBC20B2121),
        .INIT_17(256'hC6A0C18F3C0DFCC338AB32AF155BCAE50AFB210977CDF5D1C11FB7790AE409CB),
        .INIT_18(256'h7C4F937D0994C3C10B21CD2F7A4F2F7B0682CD0975CD0988CD5A1614F6C39FFF),
        .INIT_19(256'h03C4C30FF70B22C3AF4738003A031838463A14FBC390067338AB21001E50419A),
        .INIT_1A(256'h2B0697C2B77A067ECD0972CDD703DBC3161EC0E1B57C23384D2AE503C4C310F7),
        .INIT_1B(256'hCDC912D10B54CD2CCFD50B88CD0682CD0972CD0B36C31A0B88CD0682CDC97BD7),
        .INIT_1C(256'hF8182B0BC8027EE7C1E3C50BA9CDC90697D2E1E72FFF21E5C9E10682CDE50985),
        .INIT_1D(256'h0CF7C003DBC3000C11D8E1390338679CFF3E6F95D03EE53E0909000638DA2AE5),
        .INIT_1E(256'h2238D62A0C05CDAF38C12238AD2A38CE222B384F2A38D62223772377AF384F2A),
        .INIT_1F(256'hE538DE2238CB3238D422676FAF19BECD38AF221FD8CDF9384B2AC138DA2238D8),
        .INIT_20(256'hC0C9EB38DC222B06F3D2D16960049FCDE5069CCDEB0E28384F2AEBC938CE2AC5),
        .INIT_21(256'hDECD19BECD38D42238CE2A38D22209283CA47DF5384D2AC1FFF62138CE22C0F6),
        .INIT_22(256'hC3C9384D53ED38D25BED03DBCA002011B57C38D42A0402C303F4C2037321F119),
        .INIT_23(256'h12282306C5F5E5F10975CD38CB320697C210D1CD38CB32013ED7F5B7AF3E0697),
        .INIT_24(256'hF820B81B4DCD060E1BCECD1B2ECD11181B87CD1B87CD1B87CD781BBCCD1B7FCD),
        .INIT_25(256'h1CC2F1F01823771B4DCC1B8AC47EF5F10D28E723090900064EEB19EBE1F7200D),
        .INIT_26(256'h2CCFE10E2838AD2AE5D72B067BCD0BCFCA0BF7C93F5BFED841FE7E1B7EC3E11C),
        .INIT_27(256'h0BB7D2E70900280138D62AE50BB7DA579A7C5F937DEBE303C4C2D72B067BCDD5),
        .INIT_28(256'hC2039FCD38CE2210D1C4000011C9579A7C5F937D0BCFC3E138AD22E1384B22EB),
        .INIT_29(256'hCD90C1E1155BCDE51531CDE1153ACDE11253CDE5E31520CDD523F57ED5F903CA),
        .INIT_2A(256'h203EDF3F3E0D16CDD7062CC22CFE7E38CE2AF90628C36069384D22EB09281531),
        .INIT_2B(256'h20DF2B051218DF7E09282B0504DF1328050520384A325C3EB7384A3A0D85C3DF),
        .INIT_2C(256'hAFDF5C3E0728B7384A3ACE287FFE4F19DACD384A32AF010638602119EACDDF0D),
        .INIT_2D(256'h08FE00000000000D82CA15FE19E5CA0DFEC83719EACC03FE412807FE79384A32),
        .INIT_2E(256'hD1E10E9DCD38602119EACD0036E5D5C5142012FE0D81C3233E052018FE0D7CCA),
        .INIT_2F(256'h0FC9CDD50D8EC3DF042338CC3271790DF8D2073E49FE780D8EDA20FE0D8EC3C1),
        .INIT_30(256'h0A1D15D03CBBAFD801D67AC8B27BE157F11531CD0FCDCDF5C5D146234E23237E),
        .INIT_31(256'h0EB3CDE523237EC5101D010FC9CD0E5FCD1680CD0975CD14F1C33FED2823BE03),
        .INIT_32(256'h2BC9E1722373232377E538BD210EB3CD013EC9D10FBDCD6FE50E53CD46234EE1),
        .INIT_33(256'hBD110E53CD79EB23E3066BCC22FEF420B80328BA0628B70C7E23FF0EE5502206),
        .INIT_34(256'h0E5FCD2303DBC3001E11C07EE138AF22E7153DCD38AB32013E38E42238AF2A38),
        .INIT_35(256'h4F2F38C12AEB384B2AF5F10EB7F4180319F0CC0DFEDF0AC81D1C1531CD0FC9CD),
        .INIT_36(256'hC12238AD2AC50EB501F5BF03DBCA001A11F1C9F1EB2338C1220738E72309FF06),
        .INIT_37(256'h28E738D85BED38D62A0F32C20EEC01E738AF5BED38B121E538DA2AE500002138),
        .INIT_38(256'h38C5220F0AF2B709E57A1531CD0F57CAE738DA5BEDC1F0180F35CDB7237E230A),
        .INIT_39(256'h44C8B7F02356235E23237E80F6C50F2701DC28E7EB38C52AEB23090900064EE1),
        .INIT_3A(256'h4E2B462BC8B57CE1D1C9C5D5E5F1F1C1D06960E5E3E7E3E1D86960E738C12A4D),
        .INIT_3B(256'hE42AE5C50EDEC32B6960702371E10B95CD38C12A4D442B59500900266E2B2BE5),
        .INIT_3C(256'hCCCDE30FCDCDD10E50CD03DBDA001C1186E538E42AE57E0976CDE309FDCDE338),
        .INIT_3D(256'hC82D2C6F46234E23237EE3E10E7EC3E5E30991210FB4CD0FB4CDEB38BF2AE50F),
        .INIT_3E(256'h2209470520E738C12A4E1B5950D5C0EB0FE4CDEB38E42A0976CDF8181303120A),
        .INIT_3F(256'h7E38AB3257AF0FC6CDC50B3601C938AF22C0E72B2B4E2B462B38AF2AC9E138C1)
    ) ram_01(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_01), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_02;
    RAMB16_S9_S9 #(
        .INIT_00(256'h7EC3C17338BF2A0B57CD0E4ECDC91A56235E23230697CA0FF7CDC50B3601C9B7),
        .INIT_01(256'h090006686623462323E5E1C10EB3CDC5000E11780238B87EE54FE3AF10A0CD0E),
        .INIT_02(256'h050410A3CD7EEBCC18901AD5D110A0CD0E7EC30FCDCDD10FBDCD6F0E53CD4D44),
        .INIT_03(256'hBB917E4FD00006BE3DC5102701E3F129CF0B54CD2CCF052829FEFF1EC50697CA),
        .INIT_04(256'hC970E1C115E5CDD72BC5E3724619E56F66237E23235F12C3CA0FF7CDC943D847),
        .INIT_05(256'h4B5BED0EDBCD0FC9CD0B1CCAB738AB3A39000021EB38DA2AC943C5D1C129CFEB),
        .INIT_06(256'hAB3247AF03C4DA0CC5CD4E38AA32AFF6C510C7012CCFC8D72B0B1CC338C12A38),
        .INIT_07(256'hCB3AD747800F38AB323C082024D6F8300CC6CDFD38D74709380CC6CD0538D738),
        .INIT_08(256'h2A141ACA38E011E738DE2A5950E538CB32AF117ACA28D67E110EF211A0CA3D38),
        .INIT_09(256'hD5E3E11126C323232323116CCA2396781132C2239679113DCAE738D62AEB38D8),
        .INIT_0A(256'hD822696038DA22E10B92CDE5C109E538DA2A000601C5E5E3116FCAD1E70A5111),
        .INIT_0B(256'h57E338AA2AE5C9E138E422036D2138E732C9E1EB23722373D1FA20E700362B38),
        .INIT_0C(256'h11D5001E38AA22E138D02229CF1180CA2CFE7E573CEBE5E3EBF1C1067ACDC5D5),
        .INIT_0D(256'hB738AA3AEA202356235E23B87E0220B9237E2528E738DA5BED193E38D82AF5E5),
        .INIT_0E(256'hCD4F237023710697CAF100041103DBC3001011122BCA96141ACA4D44F103CDC2),
        .INIT_0F(256'hE1EB15CACDE5237023F57103C10230000B01791738AA3A237138C32223230BA0),
        .INIT_10(256'h29EB5E38C32A5703FA20E700362B38DA220BA9CD0BB7DA19EB4B42F5EA203DF1),
        .INIT_11(256'hD115CACDE511CDD2E7F5E32356235EE116237E4F472138F1237223732B2BEB09),
        .INIT_12(256'h0BCDD1C1211531CD09181531CD175721C938D02AEB09C12929E9204D443DF119),
        .INIT_13(256'h46CDF5D019FED1C11523CDEB1513CDEB3C2F0C30901523CAB738E73AC8B77815),
        .INIT_14(256'hAF52181352CD012E03D3CA34235E301310CD129FF238E421B77C1330CDF16715),
        .INIT_15(256'hFE08D6786F65544A2720B77947AF6368131CDC4F997E23579A7E235F9B7E4790),
        .INIT_16(256'hF24F8F7957177A29050B184F1F04FC301705790A20B2B57CC938E732AFF020E0),
        .INIT_17(256'h4FA980E67E23461303FCB738E72178D228D430778638E7210928B7455C7812C8),
        .INIT_18(256'h7E38E821C94F897E23578A7E235F837E03D3C3C034800EC00CC014C01C1523C3),
        .INIT_19(256'h6F09C6F518000E515A43073808D60006C94F997D579A7D5F9B7D47906FAF772F),
        .INIT_1A(256'h00EF18471F785F1F7B571F7A4F1F79C82DAF0618FA304F1FC82D790920B0B37A),
        .INIT_1B(256'h11720A834DB0E2810000000482837FA9848DCD75834363248319F79A04810000),
        .INIT_1C(256'hCDF5A838E732803E152ECD36187218118031011395CD0697EAB7EF7F3504F483),
        .INIT_1D(256'h1513CDF1142FCDD1C11846CD1374211523CDEB1513CDE1C11846CD1363211513),
        .INIT_1E(256'h21585000000138F722EB38F6327914ACCD002EC8EFD1C1211261C3D1C114F6CD),
        .INIT_1F(256'h3AE1EB1938F72AE50B3079671F082EE52C28B7237E38E421E5E513EB21E512B0),
        .INIT_20(256'h4F515A43C9E1D9207C2D4720F678042810E6471F785F1F7B571F7A4F1F8938F6),
        .INIT_21(256'h03D3CA3403D3CA3414ACCDFF2E03C7CAEFD1C11523CD0000118420011513CDC9),
        .INIT_22(256'h00DE3810CD7DC5E5381C325F574FAFEB413811327E2B3815327E2B3819327E2B),
        .INIT_23(256'h0228B5B478F5C0E61F381C3A171487F21F3D3C79E1C1D237F1F1381C3207303F),
        .INIT_24(256'h20B3B279381C3217381C3A471778294F177957177A5F177B1712F2C3B4E1203E),
        .INIT_25(256'h7780C614CCF278A81F4780AE38E7217D1D28B77812C3C3AF20E13538E721E5B7),
        .INIT_26(256'h4703D3DA02C6C8B778152ECD03D3C312C3F2E1B7E12FEFC92B771546CD141ACA),
        .INIT_27(256'h704F38E7210000118806EFC93CC09F172FFE38E63A03D3C3C03438E7211261CD),
        .INIT_28(256'hC9EBE5E338E62AE5E338E42AEBC97780EE7E38E621F0EF12ADC3178036230006),
        .INIT_29(256'h1A040638E411C92346234E2356235E38E421C9EB38E622696038E422EB1531CD),
        .INIT_2A(256'h0028CAB778C9AE1F4F1F3707797723231F3F771F37077E38E621C9FA10231377),
        .INIT_2B(256'h2BC0BE7A2BC0BE792BC0BE7823C9A91F1573CDF879AE38E621C879EFE514EF21),
        .INIT_2C(256'h177C1330CD90983E15AAFC67AE1546CD152ECDE5C8B75F574F47C9E1E1C0967B),
        .INIT_2D(256'h361586CD7ED038E43A98FE7E38E721C90BC03CA37A1BC9E1131CDC00061303DC),
        .INIT_2E(256'h11CDDA0915E0D2EB29EB11CDDA29103EC8B178000021C9F112ADCD1779F57B98),
        .INIT_2F(256'h161ACA2EFE163FDAD74F2F5F574712C3CD2B01282BFE0528F52DFEC915D2C23D),
        .INIT_30(256'h7BE515F7CA0C0C5F93AF161EC2141661DAD70A98CDD7161EC245FE160ACA65FE),
        .INIT_31(256'hD5C93DF114D4CDF5C8C9EB150BCCF1D11621C23CF11421CDF5162DF21637F490),
        .INIT_32(256'h61C3D1C114F6CD1513CD15F7C3D1C1E11656CD30D6F114D4CDD5E5C547897857),
        .INIT_33(256'h14FBCD9806AFEBD50E9C11E10E9DCD036921E5160EC35F30D686078307077B12),
        .INIT_34(256'hF8119143011748CDF5AF150BFCE51742CA3036232D36168CF22036EFE538E921),
        .INIT_35(256'h1586CD3C1250CD1748CDF53CF11421CD169BC3F51638CDF116B9E2B7155BCD4F),
        .INIT_36(256'h16E6C205175E11F5E13D3D023E473C16D5D208FE16D5FA3C81F10306011523CD),
        .INIT_37(256'h9E7923579E7A235F967B042F06E1152ECDD5E5C51538CC2E3605233036232E36),
        .INIT_38(256'h1ACA30FE7E2B1726CA0516E6C20DC12370E1EB1523CD231310CD16F5D22B2B4F),
        .INIT_39(256'h3AC61738D20AD6042F063C2F2D361736F22B362345361745CAF11538C42EFE17),
        .INIT_3A(256'h86A00F424080000000E916B0E2E1B7155BCD23F711947401C9E1712377237023),
        .INIT_3B(256'hD1C11520CD1757211513CDE9E3150B2100000100000A0000640003E800271001),
        .INIT_3C(256'hFE38E73AF517B5F2152ECD7FF679C5D512C4CAB703C7CAB7178CF217CDCA78EF),
        .INIT_3D(256'h1770DC38E422E138E622E11F7CE1155BCDF5D1C115B1CDC5D5F10F18F1033899),
        .INIT_3E(256'h3868FE223088FE38E73A13CBCDAA3B1181380113CBCDD1C11385CDC5D5150BCC),
        .INIT_3F(256'hCD13CBC34A000011C11846CD181A21125ECDF51528D1C181C615B1CD1513CD30)
    ) ram_02(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_02), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_03;
    RAMB16_S9_S9 #(
        .INIT_00(256'hE07459887C071523C300001181000103D3C312C3C3F1F1180EF2B738E63A1513),
        .INIT_01(256'hCDE5D513C9111513CD81000000803172187E75FE1A7C63505E7A1E1DC4772697),
        .INIT_02(256'hE51531CDE113CBCDE5F5C5D5C83DD1C1F1061520CD237E1513CDE113CBCD152E),
        .INIT_03(256'h87872377000607E686C83820211520CD38412118C4FA382021EFE918E11261CD),
        .INIT_04(256'h1253CD094F878718C721381F328801FE000603E63C381F3A13CBCD1531CD094F),
        .INIT_05(256'h412112B0CD1C150C770420ABD67E34381E218036462B80364F4FEE597B152ECD),
        .INIT_06(256'h38E73A1253CD1953216875D1106992E9996846B168D518772B772B77153AC338),
        .INIT_07(256'hCD1513CD13CBCDF983117E2201D5150B1138E6327FE618F3F2B738E63AD877FE),
        .INIT_08(256'h118080011261CD0000117F80011935FA155BCD0000117F0001125ECDD1C115B1),
        .INIT_09(256'h3280EE1942F2F5B738E63A150BCD1261CD0000117F0001150BF4EF1261CD0000),
        .INIT_0A(256'h861ED7FB057F00000081490FDBC938E63280EE38E63AF0F11837CD195B2138E6),
        .INIT_0B(256'hCD1523CDEB1513CDE1C118DDCD1513CD83490FDB86A55DE18723345887992665),
        .INIT_0C(256'h38463ADF203E0C2009FEF5F119D6CAB738473AF50DF703C4C30EF7142DC318D7),
        .INIT_0D(256'h32AF1AE8C3F138463219C7CC84FE3C38463A0C380B280DD6F5F1C9F1F62007E6),
        .INIT_0E(256'h003AC91A2FCD1D72C3F1C9384632AF19BBCD0A3E19BBCD0D3EC8B738463A3847),
        .INIT_0F(256'h1A18CDE5D7C9384632AF0428B738473ADF0A3EDF0D3E385F2100360518C8B738),
        .INIT_10(256'hB700367E380A21E5C9E138AB32013E38E422036D211019CD5FF10E4ECDF50928),
        .INIT_11(256'h0A2003FE1E7ECDC9FB281A39CD380A32AFC013FE380A32C81A39CDC9E11A39CC),
        .INIT_12(256'h201AB708A03602281A8ECD1A7FCD08013E0218AFC9B71FCEC30BBECCB7385E3A),
        .INIT_13(256'hCFC9E10B23CDAF001602200116A61A06201A8ECD1A7FCDD7C9E177B606A62F03),
        .INIT_14(256'h38E7D1C5004F210697DAE7004721D5C5E5E3C9C129CF1AD0CD2CCFD51AD0CD28),
        .INIT_15(256'h28B71ACA11093C013029CB07F6183D3D3D19063803FE0028117B302821C1D1F5),
        .INIT_16(256'hD1E11E64CDE51A7FCDD50682C30985CD401008040201C9AEA0F67EF9183D1304),
        .INIT_17(256'hF9201D0F1B0ACDF1081E1B08CDFA2801E6FEDBD9F5F511F70A3E1AE8CD0D3EC9),
        .INIT_18(256'h33E8113028211AE1CDD5E5C9000000FD2025B126FED3003EC9F1D91B0ACD013E),
        .INIT_19(256'h7ECD0E9DCD00B5210E9DCDF51BE821C5D5E5C9E1D11AE1CDF838E7231AE8CD7E),
        .INIT_1A(256'h7DF8202515CB1B62CD0826FB381B62CDFC0ED9C9E1D1C1F119EACDF9200DFE1E),
        .INIT_1B(256'hE5C9C949FEF93018CB40ED3CF93818CB40ED3CAFFB301F78EDFB381F78EDC9D9),
        .INIT_1C(256'hCD021EFF3E1BA5CD081EF11BA5CD011EAFF5FC0ED9F51B8ACDAD181BF721C5D5),
        .INIT_1D(256'h0C06C5F5C9C9EB201DF72005FD20256541ED0406802E0238402E17C9F1D91BA5),
        .INIT_1E(256'h0528B71B4DCDF810F8203C1B4DCD0606C5F5C9F1C11B8ACDAFF9101B8ACDFF3E),
        .INIT_1F(256'h45523C207373657250000A0D3E59414C503C207373657250C9F1C1EB18F7283C),
        .INIT_20(256'hCDAF0F061D38CD384F2A1D25CDE51CB8CD0C62CAAAFE15F7000A0D3E44524F43),
        .INIT_21(256'hFF3EF501FE232F01AF022895D60C63CAAAFE14F7C9E11D4BCD1F4001FB101B8A),
        .INIT_22(256'h1D0DCD1D06211228D11CEDCD3857211CD9CD1B2ECDD5385D32AF1CB1CD385E32),
        .INIT_23(256'h5E3201FE38E43A0BBEDC38E432F11D0DCD1CFE21DA18F810F820B71B4DCD0A06),
        .INIT_24(256'hE738D62AEB230480C3385E32FF3E0E9DCD036E2138D62211201D51CD384F2A38),
        .INIT_25(256'h2B1006CDE50985CDC8D72B385132AF000A0D6461420401C30E9DCD1CAB21EA38),
        .INIT_26(256'h385D32AF1BCECDC9E1FB1023003641F71008280D1323771A385121060E462B2B),
        .INIT_27(256'h6F46C9F8201DC00323BE0AC8B70A061E385101C9F91023771B4DCD0606385721),
        .INIT_28(256'hCDF810DF0128B7237E06063857210E9DCDF5D500203A70696B5300203A646E75),
        .INIT_29(256'h1A38D62AEB1BBCCDC9F9101B8ACD237E38512106061BBCCD1B7FCDC9D1F119EA),
        .INIT_2A(256'h4DCD0A06572F9F385D32FF3E1BCECDC9FB20B1780B000001C9F820E71B8ACD13),
        .INIT_2B(256'h3A1420B738003A1A280AFEF513F7C9AFEE10EE2023B77E0BA9CD73C0A2965F1B),
        .INIT_2C(256'h1E45CA0BFE1E14CA07FED9F5F11A2FCD380832173E08203808323D0E28B73808),
        .INIT_2D(256'h5BED2C181E1FCD7738012A13280AFE0D280DFE302808FE7B77380D3A38012A5F),
        .INIT_2E(256'h38003A0D181DFECD1218380122190028111DD8D2E733C0111F1852ED57AF3800),
        .INIT_2F(256'h9801C977380D3A38012AC9F1D97F36380D327E38012A1E3ECD20363D2B0228B7),
        .INIT_30(256'h2AD4181E64CD00321100C801C9FB1023203633C1212806B0ED30502130281103),
        .INIT_31(256'h01221DFEC31E3ECD33C1210938003EE733E8112323133826FE3C2338003A3801),
        .INIT_32(256'h7A1B237003FF111DE7C3AF3029211E59CD06061E59CD3000212006C938003238),
        .INIT_33(256'h12F7FA182BC8B57CE1D5EE180B1E76CDFCD33C1E76CDFCD3AFC8B178C9F920B3),
        .INIT_34(256'h32AF1F36F2B7380B227E23EB05363C380FFE7E34380F21EB1A28B77C380B2AD9),
        .INIT_35(256'h203FE62F78EDBF061F200FE62F78ED7F061628380E213FE62F78ED00FF01380C),
        .INIT_36(256'hCB7BFC301F1C000011F71800362B34C9D9AF3404280338BE463E23F53808CB16),
        .INIT_37(256'hF9180036C9D9AF06360218340C280538BE043E0F202377BE5FF81806C6043018),
        .INIT_38(256'hF2B7007EDD19DD1F3721DD04281F6521DD67CB0C281F9321DD6FCB78ED7F0634),
        .INIT_39(256'h2F2D2E3B0D3A083DC9D97FE6380B22F7200D1F28F2B77E230244214F7FD61F36),
        .INIT_3A(256'h7A7365337864723474356663766779366268753769386A6E6D6B6F392C6C7030),
        .INIT_3B(256'h59264248552749284A4E4D4B4F293C4C503F5E5F3E400D2A5C2B713177326120),
        .INIT_3C(256'hC3CA10301E81C4940DC11C825121572241205A53452358445224542546435647),
        .INIT_3D(256'h8E979BC69A13858A188612A584888303C7071990C908158C098D9CC80D9D0F92),
        .INIT_3E(256'h38B12138F9222B2B0C20CD38CE2AF938F92A1A25C3E138F92239000421E51189),
        .INIT_3F(256'hF5F5F5F5F5F5F5F50E9DC3015F212010C3380932FFD3AA3E0041C3FED3FF3EC9)
    ) ram_03(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_03), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_04;
    RAMB16_S9_S9 #(
        .INIT_00(256'hE0D3013EF3D3133EF2D3223EF1D3213EF0D3C03E38A03120D3C3207EC32009C3),
        .INIT_01(256'h01111FE1C325EFCD013E205ECDF620150423EBD37E41ED20160006EA0E203E21),
        .INIT_02(256'hF1DB03330B2202D40FF704190C2C03BB0CCC0FFF03CC0F1F022E0FF101F10F11),
        .INIT_03(256'hFF21C9F1D3F1F2D3F1B0ED080001B00021400011F2D3003EF1D3153EF5F2DBF5),
        .INIT_04(256'h1FF2CD38062220F1210BBECD384F22230036390021384B2219FFCE1138AD22BE),
        .INIT_05(256'h0D0153C319EACD19EACDF5181D72CD0528B72602CD25EFCD023E0E9DCD20BF21),
        .INIT_06(256'h11F2D3233EE010C320DBC200FE00206D6574737953202B73756972617571410A),
        .INIT_07(256'h79B1ED000601C5211321E5237EF5E328F9C3F3D3233EB0ED400001C000218000),
        .INIT_08(256'h21A62193217F210F1B0A161718C9E3F1E1E96F66237E678CAF6F8521182187C1),
        .INIT_09(256'h4C4C41C347554245C44753D05455CF455441434FCC534CC3544944C521D421B8),
        .INIT_0A(256'hEF80245845C8594FCA4EC944C34C45C45249444BCD5249C4455641D344414FCC),
        .INIT_0B(256'hC122C22280226C239F238E23CD23DE2353230422FC21EF224321F4220421F021),
        .INIT_0C(256'h2311EBC5E1F1C1210FC2CBFE782105C3217921E5872FD6D032FED82FFEC5E1F1),
        .INIT_0D(256'hD6C9C50230E1F1C105A8C32124114FD3D6C9D50230D4FEE1F1D104F9C3D30621),
        .INIT_0E(256'h3AE10985CDE50BCBCAE1F1F10665C3215F21EB00064F0703C4D20DFE03C4DA54),
        .INIT_0F(256'h0B54CD2CCFD50682CD0972CDC9DF0B3EC906DBC3062C010BCFCD28A5CA3D38AB),
        .INIT_10(256'hEB2221CDEB57F11C0697D218FE0B54CD2CCF0697D226FE3DF50B54CDC979EDC1),
        .INIT_11(256'h19300011192929293D7B6F6200165AEB8587877DE177380D3A38012AD9E5F5C9),
        .INIT_12(256'hD6E91823C02CFE7EF6D30B54CD2CCFF7D3103010FE0B54CD03D6CA00FE1DE7C3),
        .INIT_13(256'h0B36C378ED4B420682CDD50A4911E30A37CD23E1EC18F8D30B54CD2CCFF9D310),
        .INIT_14(256'hED0E3E0F2843CBFF3E00F7015F033E0220B77B0682CDD50A4911E30A37CD23E1),
        .INIT_15(256'hC32FFC1078EDFF060D79ED0F3E00F7010E284BCB1220FFFEFC1078EDFF060D79),
        .INIT_16(256'h003622E6CD7B22E6CD7A0428B77A38E9210682CDD50A4911E30A37CD23E10B36),
        .INIT_17(256'hCD0972CDC9237730C607C602380AFE0FE67822EFCD1F1F1F1F470E2FC338E921),
        .INIT_18(256'hED0682CD0972CD0D28AAFE2786CD27F3C22CFE2787CD26B4CD26E8CDC9D50682),
        .INIT_19(256'h60E50975CD0697C238CB3210D1CD38CB32013E2327C5C3232CCD27B3C3BFFC53),
        .INIT_1A(256'h30C22CFE2787CD26B4CD26E8CDC9E1BFFE53ED1B1B1BBFFC2223090900064E69),
        .INIT_1B(256'h82CD0972CD2303D6C22CFE2787CDBFFC53ED0682CD0972CD2028AAFE2786CD28),
        .INIT_1C(256'hE5C9E126E0CD26D3CD25EFCD193EE526B4CD2867C3232CCD2892C3BFFE53ED06),
        .INIT_1D(256'hE526B4CDE1C9E119EACDF5181D72CD0528B72602CD26E0CD25EFCD1E3E1820B7),
        .INIT_1E(256'hB7E5C9E126E0CD26D3CD25EFCD1B3EE526B4CDEC1826E0CD26D3CD25EFCD1C3E),
        .INIT_1F(256'h183E26E0CD26D3CD25EFCD163E26E8CDE526B4CDE10518BF0132BF0032AF0920),
        .INIT_20(256'h322602CD2557C3E1241CF2B72545CAFCFE2602CD260BCDAF25EFCD183E380832),
        .INIT_21(256'h3FCB3FCB1F38523A1F38533A1D72CD2D3E2616CD50C63FCB3853322602CD3852),
        .INIT_22(256'hCD3852322602CD1D72CD203E2616CD1FE638523A1D72CD2D3E2616CD3FCB3FCB),
        .INIT_23(256'hCB1F39CB38523A4F07E638533A1D72CD3A3E2616CD3FCB3FCB3FCB3853322602),
        .INIT_24(256'h02CD2602CD0E9DCD253E21142847CB2602CD2616CD1F39CB1F39CB1F39CB1F39),
        .INIT_25(256'h55322602CD3854322602CD3853322602CD3852322602CD7F182602CD2602CD26),
        .INIT_26(256'h6F38523A6738533A1220FCE638533A1920B738543A3B20F0E638543A4220B738),
        .INIT_27(256'h3E2635CD1DCB3CCB1DCB3CCB6F38533A670FE638543A3E181D72CD423E2635CD),
        .INIT_28(256'h35CD1DCB3CCB1DCB3CCB1DCB3CCB1DCB3CCB6F38543A6738553A22181D72CD4B),
        .INIT_29(256'h3C202403C319EACDF5181D72CD0528B72602CD1D72CD203E00181D72CD4D3E26),
        .INIT_2A(256'h053E023808FE3D44EDC9E12557FAB72602CD260BCDAF25EFCD173E003E524944),
        .INIT_2B(256'h25BD25AE25AA259C258E258403F4C3DF3F3E6F66237E6700CE7C6F8587257421),
        .INIT_2C(256'h61766E49006E65706F20796E616D206F6F5400646E756F6620746F4E25D325CB),
        .INIT_2D(256'h6B6E55007374736978652079646165726C4100464F45006D617261702064696C),
        .INIT_2E(256'h25E621007974706D6520746F4E006B736964206F4E00726F727265206E776F6E),
        .INIT_2F(256'hC3F1F4D3803EF618F5DB042801E6F4DBF500656C69662064614203F4C3DF3F3E),
        .INIT_30(256'h000EF81864D6043864FEC9F5D3F1FA2002E6F4DBF5C9F5DBFA2801E6F4DB260B),
        .INIT_31(256'hFC18012652CDD8F0010116C91D72CD30C6F11D72CD2FC679F50AC6FB300AD60C),
        .INIT_32(256'hC600160828B742EDFC38093CFF3EFF0E00162652CDF60E2652CDFF9C012652CD),
        .INIT_33(256'h2A38C12238AD2A38DC2238CE222B384F2AC91D72CD203EF62842CBC91D72CD30),
        .INIT_34(256'h6B62384F5BED38DE2238CB3238D422676FAF38AF2238B12138DA2238D82238D6),
        .INIT_35(256'h2323BF00320FF7CDE50985CDC9EB18722373EBFC2023BEAF2323230E28B6237E),
        .INIT_36(256'h273BC35F3CBF003A0016BF0121C9E112AFB0ED0228B74F0006BF011168662346),
        .INIT_37(256'h26E0C326D3CD260BCD003E25EFCD103E26E0C325EFCD1F3EC92557FAB72602CD),
        .INIT_38(256'h0BCD7A260BCD7B260BCDAF25EFCD123E26E0C326D3CD260BCD193E25EFCD103E),
        .INIT_39(256'h0828B37AD5C9D1F4181B23772602CD0828B37AD5572602CD5F2602CD26E0CD26),
        .INIT_3A(256'hE0CD273BCD260BCD7A260BCD7B260BCDAF25EFCD133EC9D1F4181B23260BCD7E),
        .INIT_3B(256'hCD260BCDAF260BCD7A260BCD7B260BCDAF25EFCD143EC9572602CD5F2602CD26),
        .INIT_3C(256'h0C0E25DDC20DFE7B2710CDBFEC21000D11F718C020FEC8B77E23C926E0CD260B),
        .INIT_3D(256'h2710CDFFFF11BFFC2A26F0CDE5C925DDC2B77EF6200D2325DDC2FFFE7EBFEC21),
        .INIT_3E(256'h25DDC223FE7EBFEC21060E2710CDBFEC21000611278FCD26F0CDE5C9E126E8CD),
        .INIT_3F(256'hBFEC21000611278FCD26F0CDE5C9E126E8CD2710CDBFFE5BEDBFFC2AF6200D23)
    ) ram_04(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_04), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_05;
    RAMB16_S9_S9 #(
        .INIT_00(256'h6FCD38D62223232323FB28BEAF2B26E8CD2710CDFFFF11384F2A278FCD2710CD),
        .INIT_01(256'h286121274ACD000D112823212700CDE500FFFFFFFFFFFFFFFFFFFFFFFFC9E126),
        .INIT_02(256'hE126E8CD274ACDEB52ED38D62A384F5BED274ACD000D11282321274ACD000611),
        .INIT_03(256'hBFFC2A274ACD000611288C21274ACD000D112823212700CDE5475250534142C9),
        .INIT_04(256'h274ACDBFFE5BEDBFFC2A2700CDE5232323232323C9E126E8CD274ACDBFFE5BED),
        .INIT_05(256'hCD172828C5CD28D1215FBF1603D60D3805FEBF003A26B4CD26E8CDC9E126E8CD),
        .INIT_06(256'hC00021F3D3233E26F0CD004D4F522EC9F520B7C023BE132928CD1A0BCBC327F3),
        .INIT_07(256'h860C06E00321AF26E8CDB0ED200001E00011C000210B2020FE7A2710CD400011),
        .INIT_08(256'hA33EF2D3223EF1D3213EF720B37A1B2377AE78400011C0002147AEFA20058023),
        .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC920D6D07BFED861FEE010C338A031F3D3),
        .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_24(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_26(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_27(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_29(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_2A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_2B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_2D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
    ) ram_05(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_05), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_06;
    RAMB16_S9_S9 #(
        .INIT_00(256'h00041C542C50286400041C542C504844001C08442C50484400AC60207820203C),
        .INIT_01(256'h002040FFFF402000000402FFFF0204003C4299A1A199423C000010007C001000),
        .INIT_02(256'hF0E0F0B81C0E0400002070381D0F070F183C5A181818181818181818185A3C18),
        .INIT_03(256'h30303030303CFCFCFFFFFF7E003C3C0000040E1CB8F0E0F00F070F1D38702000),
        .INIT_04(256'hDBBDFF7E003C3C003C3C3C3C3C3C3C3C0C0C0C0C0C3C3F3F0000003C3C3C3CFF),
        .INIT_05(256'hDCDF7939003C38003838181C1E1B3E7C7F7C7838003C3800C3C3C3E766663C7E),
        .INIT_06(256'h000000000F0F0F0F0F0F0F0F00000000DB99BDE724663C180080C3F33B1F3F7C),
        .INIT_07(256'hFFFFFFFF000000000F0F0F0FF0F0F0F000000000F0F0F0F0F0F0F0F000000000),
        .INIT_08(256'h0028287C287C2828000000000028282800100010101010100000000000000000),
        .INIT_09(256'h00000000001008080034485420505020000C4C20100864600010781438503C10),
        .INIT_0A(256'h000010107C101000001054381038541000100804040408100010204040402010),
        .INIT_0B(256'h00004020100804000010000000000000000000007C0000000020101000000000),
        .INIT_0C(256'h003844041808047C007C402018044438003810101010301000384464544C4438),
        .INIT_0D(256'h002020201008047C003844447840201C003844040478407C0008087C48281808),
        .INIT_0E(256'h00201010001000000000001000100000007008043C4444380038444438444438),
        .INIT_0F(256'h001000101008443800201008040810200000007C007C00000008102040201008),
        .INIT_10(256'h003844404040443800784444784444780044447C44442810003C40585C544438),
        .INIT_11(256'h003C444C4040403C004040407840407C007C40407840407C0078444444444478),
        .INIT_12(256'h004448506050484400384404040404040038101010101038004444447C444444),
        .INIT_13(256'h00384444444444380044444C546444440044444454546C44007C404040404040),
        .INIT_14(256'h0038440438404438004448507844447800344854444444380040404078444478),
        .INIT_15(256'h00446C545444444400102844444444440038444444444444001010101010107C),
        .INIT_16(256'h007C60606060607C007C40201008047C00101010102844440044442810284444),
        .INIT_17(256'h007C0000000000000000004428100000007C0C0C0C0C0C7C0000040810204000),
        .INIT_18(256'h001C2020201C0000005864446458404000344C444C3400000000000000102020),
        .INIT_19(256'h38043C444C34000000101010381010080038407C4438000000344C444C340404),
        .INIT_1A(256'h0044487050484040300808080808000800381010103000100044444444784040),
        .INIT_1B(256'h0038444444380000004444444478000000525252526C00000038101010101030),
        .INIT_1C(256'h00780438403C0000004040406058000006344C444C3400004058644464580000),
        .INIT_1D(256'h002C5252525200000010282844440000003C44444444000000101010107C1010),
        .INIT_1E(256'h000C10102010100C007C2010087C000038043C24242400000044281028440000),
        .INIT_1F(256'hFFFFFFFFFFFFFFFF000000403804000000601010081010600010101000101010),
        .INIT_20(256'h1C1C183878D87C3EFE3E1E1C003C1C008080808080808080FFFFFFFFFFFFFF00),
        .INIT_21(256'h00183C7E7E3C180055AA55AA55AA55AA50A050A050A050A055AA55AA00000000),
        .INIT_22(256'h18183C7EFFDB183C3C18DBFF7E3C1818FFFFFFFFFFFF0000FFFF000000000000),
        .INIT_23(256'hFFFF7E7E3C3C1818C0F0FCFFFFFCF0C00001C3CFDCF8FC3E3BFB9E9C003C1C00),
        .INIT_24(256'hBCBCFF3D013C4A3C3D3DFFBC803C523CFEFEFEFEFEFEFEFEFF00000000000000),
        .INIT_25(256'hC0C0C0C0C0C0C0C03C7EFFFFFFFF7E3C050A050A050A050A0000000055AA55AA),
        .INIT_26(256'h0C1C39FFFF391C0C30389CFFFF9C3830F8F8F8F8F8F8F8F8E0E0E0E0E0E0E0E0),
        .INIT_27(256'h18183C3C7E7EFFFF030F3FFFFF3F0F0300667E42C3FF18000018FFC3427E6600),
        .INIT_28(256'h0000000000FFFFFF00000000000F0F0F0000000000F0F0F00000000000000000),
        .INIT_29(256'h000000F0F0FFFFFF000000F0F00F0F0F000000F0F0F0F0F0000000F0F0000000),
        .INIT_2A(256'h0000000F0FFFFFFF0000000F0F0F0F0F0000000F0FF0F0F00000000F0F000000),
        .INIT_2B(256'h000000FFFFFFFFFF000000FFFF0F0F0F000000FFFFF0F0F0000000FFFF000000),
        .INIT_2C(256'hF0F0F00000FFFFFFF0F0F000000F0F0FF0F0F00000F0F0F0F0F0F00000000000),
        .INIT_2D(256'hF0F0F0F0F0FFFFFFF0F0F0F0F00F0F0FF0F0F0F0F0F0F0F0F0F0F0F0F0000000),
        .INIT_2E(256'hF0F0F00F0FFFFFFFF0F0F00F0F0F0F0FF0F0F00F0FF0F0F0F0F0F00F0F000000),
        .INIT_2F(256'hF0F0F0FFFFFFFFFFF0F0F0FFFF0F0F0FF0F0F0FFFFF0F0F0F0F0F0FFFF000000),
        .INIT_30(256'hFCFCFCFCFCFCFCFC000000003C7EFFFFFFFEFCF8F0E0C080FF7F3F1F0F070301),
        .INIT_31(256'h0000000003070F0F0000001818000000183C7EFFFF7E3C1800003C3C3C3C0000),
        .INIT_32(256'h03070F0F0F0F07038040201008040201F0F0E0C000000000181818FFFF181818),
        .INIT_33(256'h0000001F1F181818181818F8F80000001818181F1F181818000000FFFF181818),
        .INIT_34(256'h0004345C3A2C1000FFFF7E3C000000004A23B411C42D44520208401180042009),
        .INIT_35(256'h0F0F07030000000018181818181818183C1842E742183C1818183C7EFFFFFF66),
        .INIT_36(256'hC0E0F0F0F0F0E0C0010204081020408000000000C0E0F0F08142241818244281),
        .INIT_37(256'h000000F8F81818181818181F1F000000181818F8F8181818181818FFFF000000),
        .INIT_38(256'h0F0F0F0000FFFFFF0F0F0F00000F0F0F0F0F0F0000F0F0F00F0F0F0000000000),
        .INIT_39(256'h0F0F0FF0F0FFFFFF0F0F0FF0F00F0F0F0F0F0FF0F0F0F0F00F0F0FF0F0000000),
        .INIT_3A(256'h0F0F0F0F0FFFFFFF0F0F0F0F0F0F0F0F0F0F0F0F0FF0F0F00F0F0F0F0F000000),
        .INIT_3B(256'h0F0F0FFFFFFFFFFF0F0F0FFFFF0F0F0F0F0F0FFFFFF0F0F00F0F0FFFFF000000),
        .INIT_3C(256'hFFFFFF0000FFFFFFFFFFFF00000F0F0FFFFFFF0000F0F0F0FFFFFF0000000000),
        .INIT_3D(256'hFFFFFFF0F0FFFFFFFFFFFFF0F00F0F0FFFFFFFF0F0F0F0F0FFFFFFF0F0000000),
        .INIT_3E(256'hFFFFFF0F0FFFFFFFFFFFFF0F0F0F0F0FFFFFFF0F0FF0F0F0FFFFFF0F0F000000),
        .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0F0F0FFFFFFFFFFFF0F0F0FFFFFFFFFF000000)
    ) ram_06(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_06), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_07;
    RAMB16_S9_S9 #(
        .INIT_00(256'h00081C3E7F7F7F367EFFE7C3FFDBFF7E7E8199BD81A5817E0000000000000000),
        .INIT_01(256'h0000183C3C1800003C18DBFFFF7E3C183C18DBE7E73C3C1800081C3E7F3E1C08),
        .INIT_02(256'h78CCCCCC7D0F070FFFC399BDBD99C3FF003C664242663C00FFFFE7C3C3E7FFFF),
        .INIT_03(256'h995A3CE7E73C5A99C0E66763637F637FE0F07030303F333F187E183C6666663C),
        .INIT_04(256'h0066006666666666183C7E18187E3C1800020E3EFE3E0E020080E0F8FEF8E080),
        .INIT_05(256'hFF183C7E187E3C18007E7E7E0000000078CC386C6C38663C001B1B1B7BDBDB7F),
        .INIT_06(256'h0010307F7F30100000080CFEFE0C080000183C7E1818181800181818187E3C18),
        .INIT_07(256'h0000183C7EFFFF000000FFFF7E3C180000002466FF6624000000FEC0C0C00000),
        .INIT_08(256'h006C6CFE6CFE6C6C000000000066666600180000181818180000000000000000),
        .INIT_09(256'h00000000003018180076CCDC76386C3800466630180C666200187C063C603E18),
        .INIT_0A(256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C),
        .INIT_0B(256'h0080C06030180C060018180000000000000000007E0000003018180000000000),
        .INIT_0C(256'h003C66061C06663C007E60300C06663C007E181818381818003C6666766E663C),
        .INIT_0D(256'h001818180C06667E003C66667C60663C003C6606067C607E0006067F66361E0E),
        .INIT_0E(256'h30181800001818000018180000181800003C66063E66663C003C66663C66663C),
        .INIT_0F(256'h001800180C06663C0030180C060C18300000007E007E0000000C18306030180C),
        .INIT_10(256'h003C66606060663C007C66667C66667C006666667E663C18003C62606E6E663C),
        .INIT_11(256'h003C66666E60663C006060607860607E007E60607860607E00786C6666666C78),
        .INIT_12(256'h00666C7870786C6600386C0C0C0C0C1E003C18181818183C006666667E666666),
        .INIT_13(256'h003C66666666663C0066666E7E7E7666006363636B7F7763007E606060606060),
        .INIT_14(256'h003C66063C60663C00666C787C66667C000E3C666666663C006060607C66667C),
        .INIT_15(256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E),
        .INIT_16(256'h003C30303030303C007E6030180C067E001818183C6666660066663C183C6666),
        .INIT_17(256'h00FE00000000000000000000C66C3810003C0C0C0C0C0C3C0002060C183060C0),
        .INIT_18(256'h003C6060603C0000007C6666667C6060003E663E063C00000000000000183030),
        .INIT_19(256'h7C063E66663E0000001818183E18180E003C607E663C0000003E6666663E0606),
        .INIT_1A(256'h00666C786C6660607018181818380018003C18181838001800666666667C6060),
        .INIT_1B(256'h003C6666663C000000666666667C000000636B7F7F660000003C181818181838),
        .INIT_1C(256'h007C063C603E000000606060667C000006063E66663E000060607C66667C0000),
        .INIT_1D(256'h00363E7F6B63000000183C6666660000003E666666660000000E1818187E1818),
        .INIT_1E(256'h000E18187018180E007E30180C7E0000780C3E666666000000663C183C660000),
        .INIT_1F(256'h00FEC6C66C38100000000000DC760000007018180E1818700018181800181818),
        .INIT_20(256'h003E663E063C423C003C607E663C000E003E666666006600780C1878CCC0CC78),
        .INIT_21(256'h1C063C60603C0000003E663E063C1818003E663E063C0070003E663E063C0066),
        .INIT_22(256'h003C181838006600003C607E663C0070003C607E663C0066003C607E663CC37E),
        .INIT_23(256'h00667E663C001818006666667E663C5A003C181838001020003C181838002418),
        .INIT_24(256'h003C66663C00663C00CECCCCFECC6C3E007FCC7F0C7F0000007E6078607E001C),
        .INIT_25(256'h003E666666007000003E66666600663C003C66663C007000003C66663C006600),
        .INIT_26(256'h18187EC0C07E1818003C666666660066003C666666663CC3780C3E6666006600),
        .INIT_27(256'h70D818183C181B0EC7C6CFC6FACCCCF83030FC30FC78CCCC00FC62307C30120C),
        .INIT_28(256'h003E666666000E00003C66663C000E00003C181838001008003E663E063C000E),
        .INIT_29(256'h00007C00386C6C3800007E003E6C6C3C00666E7E7666007E006666667C007C00),
        .INIT_2A(256'h0FCC6633DECCC6C3000006067E000000000060607E000000003C666030180018),
        .INIT_2B(256'h0000CC663366CC0000003366CC663300001818181800181803CF6F37DBCCC6C3),
        .INIT_2C(256'h1818181818181818EEBBEEBBEEBBEEBBAA55AA55AA55AA558822882288228822),
        .INIT_2D(256'h363636FE00000000363636F636363636181818F818F81818181818F818181818),
        .INIT_2E(256'h363636F606FE00003636363636363636363636F606F63636181818F818F80000),
        .INIT_2F(256'h181818F800000000000000F818F81818000000FE36363636000000FE06F63636),
        .INIT_30(256'h1818181F18181818181818FF00000000000000FF181818180000001F18181818),
        .INIT_31(256'h36363637363636361818181F181F1818181818FF18181818000000FF00000000),
        .INIT_32(256'h363636F700FF0000000000FF00F7363636363637303F00000000003F30373636),
        .INIT_33(256'h000000FF00FF1818363636F700F73636000000FF00FF00003636363730373636),
        .INIT_34(256'h0000003F36363636363636FF00000000181818FF00FF0000000000FF36363636),
        .INIT_35(256'h363636FF363636363636363F000000001818181F181F00000000001F181F1818),
        .INIT_36(256'hFFFFFFFFFFFFFFFF1818181F00000000000000F818181818181818FF18FF1818),
        .INIT_37(256'h00000000FFFFFFFF0F0F0F0F0F0F0F0FF0F0F0F0F0F0F0F0FFFFFFFF00000000),
        .INIT_38(256'h0036363636367F00006060606060667E006663636C66663C003B6E646E3B0000),
        .INIT_39(256'h000C0C0C0C6E3B0060303E333333330000386C6C6C3F0000007E66301830667E),
        .INIT_3A(256'h003C66663E0C180E007736366363361C001C36637F63361C7E183C66663C187E),
        .INIT_3B(256'h006666666666663C001C30607C60301CC0607EDBDB7E0C0600007EDBDB7E0000),
        .INIT_3C(256'h007E000C1830180C007E0030180C1830007E0018187E181800007E007E007E00),
        .INIT_3D(256'h0000DC7600DC7600001818007E00181870D8D8181818181818181818181B1B0E),
        .INIT_3E(256'h1C3C6CEC0C0C0C0F0000001800000000000000181800000000000000386C6C38),
        .INIT_3F(256'h000000000000000000003C3C3C3C00000000003C30180C380000006C6C6C6C78)
    ) ram_07(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_07), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_08;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_08(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_08), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_09;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_09(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_09), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_10;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_10(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_10), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_11;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_11(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_11), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_12;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_12(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_12), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_13;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_13(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_13), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_14;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_14(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_14), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_15;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_15(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_15), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_16;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_16(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_16), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_17;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_17(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_17), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_18;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_18(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_18), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    wire [7:0] rddata_19;
    RAMB16_S9_S9 #(
        .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram_19(
        .CLKA(clk), .SSRA(1'b0), .ADDRA(addr[10:0]), .DOA(rddata_19), .DOPA(), .DIA(8'b0), .DIPA(1'b0), .ENA(1'b1), .WEA(1'b0),
        .CLKB(clk), .SSRB(1'b0), .ADDRB(11'b0),      .DOB(),          .DOPB(), .DIB(8'b0), .DIPB(1'b0), .ENB(1'b1), .WEB(1'b0));

    always @* case (addr[15:11])
        5'd0: rddata <= rddata_00;
        5'd1: rddata <= rddata_01;
        5'd2: rddata <= rddata_02;
        5'd3: rddata <= rddata_03;
        5'd4: rddata <= rddata_04;
        5'd5: rddata <= rddata_05;
        5'd6: rddata <= rddata_06;
        5'd7: rddata <= rddata_07;
        5'd8: rddata <= rddata_08;
        5'd9: rddata <= rddata_09;
        5'd10: rddata <= rddata_10;
        5'd11: rddata <= rddata_11;
        5'd12: rddata <= rddata_12;
        5'd13: rddata <= rddata_13;
        5'd14: rddata <= rddata_14;
        5'd15: rddata <= rddata_15;
        5'd16: rddata <= rddata_16;
        5'd17: rddata <= rddata_17;
        5'd18: rddata <= rddata_18;
        5'd19: rddata <= rddata_19;
        default: rddata <= 8'h00;
    endcase

endmodule
