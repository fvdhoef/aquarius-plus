module charram(
    input  wire        clk,

    // input  wire [10:0] addr1,
    // output reg   [7:0] rddata1,
    // input  wire  [7:0] wrdata1,
    // input  wire        wren1,

    input  wire [10:0] addr2,
    output reg   [7:0] rddata2);

    reg [7:0] ram [2047:0];

    initial begin
        ram[   0] = 8'h3C; ram[   1] = 8'h20; ram[   2] = 8'h20; ram[   3] = 8'h78;
        ram[   4] = 8'h20; ram[   5] = 8'h60; ram[   6] = 8'hAC; ram[   7] = 8'h00;
        ram[   8] = 8'h44; ram[   9] = 8'h48; ram[  10] = 8'h50; ram[  11] = 8'h2C;
        ram[  12] = 8'h44; ram[  13] = 8'h08; ram[  14] = 8'h1C; ram[  15] = 8'h00;
        ram[  16] = 8'h44; ram[  17] = 8'h48; ram[  18] = 8'h50; ram[  19] = 8'h2C;
        ram[  20] = 8'h54; ram[  21] = 8'h1C; ram[  22] = 8'h04; ram[  23] = 8'h00;
        ram[  24] = 8'h64; ram[  25] = 8'h28; ram[  26] = 8'h50; ram[  27] = 8'h2C;
        ram[  28] = 8'h54; ram[  29] = 8'h1C; ram[  30] = 8'h04; ram[  31] = 8'h00;
        ram[  32] = 8'h00; ram[  33] = 8'h10; ram[  34] = 8'h00; ram[  35] = 8'h7C;
        ram[  36] = 8'h00; ram[  37] = 8'h10; ram[  38] = 8'h00; ram[  39] = 8'h00;
        ram[  40] = 8'h3C; ram[  41] = 8'h42; ram[  42] = 8'h99; ram[  43] = 8'hA1;
        ram[  44] = 8'hA1; ram[  45] = 8'h99; ram[  46] = 8'h42; ram[  47] = 8'h3C;
        ram[  48] = 8'h00; ram[  49] = 8'h04; ram[  50] = 8'h02; ram[  51] = 8'hFF;
        ram[  52] = 8'hFF; ram[  53] = 8'h02; ram[  54] = 8'h04; ram[  55] = 8'h00;
        ram[  56] = 8'h00; ram[  57] = 8'h20; ram[  58] = 8'h40; ram[  59] = 8'hFF;
        ram[  60] = 8'hFF; ram[  61] = 8'h40; ram[  62] = 8'h20; ram[  63] = 8'h00;
        ram[  64] = 8'h18; ram[  65] = 8'h3C; ram[  66] = 8'h5A; ram[  67] = 8'h18;
        ram[  68] = 8'h18; ram[  69] = 8'h18; ram[  70] = 8'h18; ram[  71] = 8'h18;
        ram[  72] = 8'h18; ram[  73] = 8'h18; ram[  74] = 8'h18; ram[  75] = 8'h18;
        ram[  76] = 8'h18; ram[  77] = 8'h5A; ram[  78] = 8'h3C; ram[  79] = 8'h18;
        ram[  80] = 8'h0F; ram[  81] = 8'h07; ram[  82] = 8'h0F; ram[  83] = 8'h1D;
        ram[  84] = 8'h38; ram[  85] = 8'h70; ram[  86] = 8'h20; ram[  87] = 8'h00;
        ram[  88] = 8'h00; ram[  89] = 8'h04; ram[  90] = 8'h0E; ram[  91] = 8'h1C;
        ram[  92] = 8'hB8; ram[  93] = 8'hF0; ram[  94] = 8'hE0; ram[  95] = 8'hF0;
        ram[  96] = 8'h00; ram[  97] = 8'h20; ram[  98] = 8'h70; ram[  99] = 8'h38;
        ram[ 100] = 8'h1D; ram[ 101] = 8'h0F; ram[ 102] = 8'h07; ram[ 103] = 8'h0F;
        ram[ 104] = 8'hF0; ram[ 105] = 8'hE0; ram[ 106] = 8'hF0; ram[ 107] = 8'hB8;
        ram[ 108] = 8'h1C; ram[ 109] = 8'h0E; ram[ 110] = 8'h04; ram[ 111] = 8'h00;
        ram[ 112] = 8'h00; ram[ 113] = 8'h3C; ram[ 114] = 8'h3C; ram[ 115] = 8'h00;
        ram[ 116] = 8'h7E; ram[ 117] = 8'hFF; ram[ 118] = 8'hFF; ram[ 119] = 8'hFF;
        ram[ 120] = 8'hFC; ram[ 121] = 8'hFC; ram[ 122] = 8'h3C; ram[ 123] = 8'h30;
        ram[ 124] = 8'h30; ram[ 125] = 8'h30; ram[ 126] = 8'h30; ram[ 127] = 8'h30;
        ram[ 128] = 8'hFF; ram[ 129] = 8'h3C; ram[ 130] = 8'h3C; ram[ 131] = 8'h3C;
        ram[ 132] = 8'h3C; ram[ 133] = 8'h00; ram[ 134] = 8'h00; ram[ 135] = 8'h00;
        ram[ 136] = 8'h3F; ram[ 137] = 8'h3F; ram[ 138] = 8'h3C; ram[ 139] = 8'h0C;
        ram[ 140] = 8'h0C; ram[ 141] = 8'h0C; ram[ 142] = 8'h0C; ram[ 143] = 8'h0C;
        ram[ 144] = 8'h3C; ram[ 145] = 8'h3C; ram[ 146] = 8'h3C; ram[ 147] = 8'h3C;
        ram[ 148] = 8'h3C; ram[ 149] = 8'h3C; ram[ 150] = 8'h3C; ram[ 151] = 8'h3C;
        ram[ 152] = 8'h00; ram[ 153] = 8'h3C; ram[ 154] = 8'h3C; ram[ 155] = 8'h00;
        ram[ 156] = 8'h7E; ram[ 157] = 8'hFF; ram[ 158] = 8'hBD; ram[ 159] = 8'hDB;
        ram[ 160] = 8'h7E; ram[ 161] = 8'h3C; ram[ 162] = 8'h66; ram[ 163] = 8'h66;
        ram[ 164] = 8'hE7; ram[ 165] = 8'hC3; ram[ 166] = 8'hC3; ram[ 167] = 8'hC3;
        ram[ 168] = 8'h00; ram[ 169] = 8'h38; ram[ 170] = 8'h3C; ram[ 171] = 8'h00;
        ram[ 172] = 8'h38; ram[ 173] = 8'h78; ram[ 174] = 8'h7C; ram[ 175] = 8'h7F;
        ram[ 176] = 8'h7C; ram[ 177] = 8'h3E; ram[ 178] = 8'h1B; ram[ 179] = 8'h1E;
        ram[ 180] = 8'h1C; ram[ 181] = 8'h18; ram[ 182] = 8'h38; ram[ 183] = 8'h38;
        ram[ 184] = 8'h00; ram[ 185] = 8'h38; ram[ 186] = 8'h3C; ram[ 187] = 8'h00;
        ram[ 188] = 8'h39; ram[ 189] = 8'h79; ram[ 190] = 8'hDF; ram[ 191] = 8'hDC;
        ram[ 192] = 8'h7C; ram[ 193] = 8'h3F; ram[ 194] = 8'h1F; ram[ 195] = 8'h3B;
        ram[ 196] = 8'hF3; ram[ 197] = 8'hC3; ram[ 198] = 8'h80; ram[ 199] = 8'h00;
        ram[ 200] = 8'h18; ram[ 201] = 8'h3C; ram[ 202] = 8'h66; ram[ 203] = 8'h24;
        ram[ 204] = 8'hE7; ram[ 205] = 8'hBD; ram[ 206] = 8'h99; ram[ 207] = 8'hDB;
        ram[ 208] = 8'h00; ram[ 209] = 8'h00; ram[ 210] = 8'h00; ram[ 211] = 8'h00;
        ram[ 212] = 8'h0F; ram[ 213] = 8'h0F; ram[ 214] = 8'h0F; ram[ 215] = 8'h0F;
        ram[ 216] = 8'h0F; ram[ 217] = 8'h0F; ram[ 218] = 8'h0F; ram[ 219] = 8'h0F;
        ram[ 220] = 8'h00; ram[ 221] = 8'h00; ram[ 222] = 8'h00; ram[ 223] = 8'h00;
        ram[ 224] = 8'h00; ram[ 225] = 8'h00; ram[ 226] = 8'h00; ram[ 227] = 8'h00;
        ram[ 228] = 8'hF0; ram[ 229] = 8'hF0; ram[ 230] = 8'hF0; ram[ 231] = 8'hF0;
        ram[ 232] = 8'hF0; ram[ 233] = 8'hF0; ram[ 234] = 8'hF0; ram[ 235] = 8'hF0;
        ram[ 236] = 8'h00; ram[ 237] = 8'h00; ram[ 238] = 8'h00; ram[ 239] = 8'h00;
        ram[ 240] = 8'hF0; ram[ 241] = 8'hF0; ram[ 242] = 8'hF0; ram[ 243] = 8'hF0;
        ram[ 244] = 8'h0F; ram[ 245] = 8'h0F; ram[ 246] = 8'h0F; ram[ 247] = 8'h0F;
        ram[ 248] = 8'h00; ram[ 249] = 8'h00; ram[ 250] = 8'h00; ram[ 251] = 8'h00;
        ram[ 252] = 8'hFF; ram[ 253] = 8'hFF; ram[ 254] = 8'hFF; ram[ 255] = 8'hFF;
        ram[ 256] = 8'h00; ram[ 257] = 8'h00; ram[ 258] = 8'h00; ram[ 259] = 8'h00;
        ram[ 260] = 8'h00; ram[ 261] = 8'h00; ram[ 262] = 8'h00; ram[ 263] = 8'h00;
        ram[ 264] = 8'h10; ram[ 265] = 8'h10; ram[ 266] = 8'h10; ram[ 267] = 8'h10;
        ram[ 268] = 8'h10; ram[ 269] = 8'h00; ram[ 270] = 8'h10; ram[ 271] = 8'h00;
        ram[ 272] = 8'h28; ram[ 273] = 8'h28; ram[ 274] = 8'h28; ram[ 275] = 8'h00;
        ram[ 276] = 8'h00; ram[ 277] = 8'h00; ram[ 278] = 8'h00; ram[ 279] = 8'h00;
        ram[ 280] = 8'h28; ram[ 281] = 8'h28; ram[ 282] = 8'h7C; ram[ 283] = 8'h28;
        ram[ 284] = 8'h7C; ram[ 285] = 8'h28; ram[ 286] = 8'h28; ram[ 287] = 8'h00;
        ram[ 288] = 8'h10; ram[ 289] = 8'h3C; ram[ 290] = 8'h50; ram[ 291] = 8'h38;
        ram[ 292] = 8'h14; ram[ 293] = 8'h78; ram[ 294] = 8'h10; ram[ 295] = 8'h00;
        ram[ 296] = 8'h60; ram[ 297] = 8'h64; ram[ 298] = 8'h08; ram[ 299] = 8'h10;
        ram[ 300] = 8'h20; ram[ 301] = 8'h4C; ram[ 302] = 8'h0C; ram[ 303] = 8'h00;
        ram[ 304] = 8'h20; ram[ 305] = 8'h50; ram[ 306] = 8'h50; ram[ 307] = 8'h20;
        ram[ 308] = 8'h54; ram[ 309] = 8'h48; ram[ 310] = 8'h34; ram[ 311] = 8'h00;
        ram[ 312] = 8'h08; ram[ 313] = 8'h08; ram[ 314] = 8'h10; ram[ 315] = 8'h00;
        ram[ 316] = 8'h00; ram[ 317] = 8'h00; ram[ 318] = 8'h00; ram[ 319] = 8'h00;
        ram[ 320] = 8'h10; ram[ 321] = 8'h20; ram[ 322] = 8'h40; ram[ 323] = 8'h40;
        ram[ 324] = 8'h40; ram[ 325] = 8'h20; ram[ 326] = 8'h10; ram[ 327] = 8'h00;
        ram[ 328] = 8'h10; ram[ 329] = 8'h08; ram[ 330] = 8'h04; ram[ 331] = 8'h04;
        ram[ 332] = 8'h04; ram[ 333] = 8'h08; ram[ 334] = 8'h10; ram[ 335] = 8'h00;
        ram[ 336] = 8'h10; ram[ 337] = 8'h54; ram[ 338] = 8'h38; ram[ 339] = 8'h10;
        ram[ 340] = 8'h38; ram[ 341] = 8'h54; ram[ 342] = 8'h10; ram[ 343] = 8'h00;
        ram[ 344] = 8'h00; ram[ 345] = 8'h10; ram[ 346] = 8'h10; ram[ 347] = 8'h7C;
        ram[ 348] = 8'h10; ram[ 349] = 8'h10; ram[ 350] = 8'h00; ram[ 351] = 8'h00;
        ram[ 352] = 8'h00; ram[ 353] = 8'h00; ram[ 354] = 8'h00; ram[ 355] = 8'h00;
        ram[ 356] = 8'h10; ram[ 357] = 8'h10; ram[ 358] = 8'h20; ram[ 359] = 8'h00;
        ram[ 360] = 8'h00; ram[ 361] = 8'h00; ram[ 362] = 8'h00; ram[ 363] = 8'h7C;
        ram[ 364] = 8'h00; ram[ 365] = 8'h00; ram[ 366] = 8'h00; ram[ 367] = 8'h00;
        ram[ 368] = 8'h00; ram[ 369] = 8'h00; ram[ 370] = 8'h00; ram[ 371] = 8'h00;
        ram[ 372] = 8'h00; ram[ 373] = 8'h00; ram[ 374] = 8'h10; ram[ 375] = 8'h00;
        ram[ 376] = 8'h00; ram[ 377] = 8'h04; ram[ 378] = 8'h08; ram[ 379] = 8'h10;
        ram[ 380] = 8'h20; ram[ 381] = 8'h40; ram[ 382] = 8'h00; ram[ 383] = 8'h00;
        ram[ 384] = 8'h38; ram[ 385] = 8'h44; ram[ 386] = 8'h4C; ram[ 387] = 8'h54;
        ram[ 388] = 8'h64; ram[ 389] = 8'h44; ram[ 390] = 8'h38; ram[ 391] = 8'h00;
        ram[ 392] = 8'h10; ram[ 393] = 8'h30; ram[ 394] = 8'h10; ram[ 395] = 8'h10;
        ram[ 396] = 8'h10; ram[ 397] = 8'h10; ram[ 398] = 8'h38; ram[ 399] = 8'h00;
        ram[ 400] = 8'h38; ram[ 401] = 8'h44; ram[ 402] = 8'h04; ram[ 403] = 8'h18;
        ram[ 404] = 8'h20; ram[ 405] = 8'h40; ram[ 406] = 8'h7C; ram[ 407] = 8'h00;
        ram[ 408] = 8'h7C; ram[ 409] = 8'h04; ram[ 410] = 8'h08; ram[ 411] = 8'h18;
        ram[ 412] = 8'h04; ram[ 413] = 8'h44; ram[ 414] = 8'h38; ram[ 415] = 8'h00;
        ram[ 416] = 8'h08; ram[ 417] = 8'h18; ram[ 418] = 8'h28; ram[ 419] = 8'h48;
        ram[ 420] = 8'h7C; ram[ 421] = 8'h08; ram[ 422] = 8'h08; ram[ 423] = 8'h00;
        ram[ 424] = 8'h7C; ram[ 425] = 8'h40; ram[ 426] = 8'h78; ram[ 427] = 8'h04;
        ram[ 428] = 8'h04; ram[ 429] = 8'h44; ram[ 430] = 8'h38; ram[ 431] = 8'h00;
        ram[ 432] = 8'h1C; ram[ 433] = 8'h20; ram[ 434] = 8'h40; ram[ 435] = 8'h78;
        ram[ 436] = 8'h44; ram[ 437] = 8'h44; ram[ 438] = 8'h38; ram[ 439] = 8'h00;
        ram[ 440] = 8'h7C; ram[ 441] = 8'h04; ram[ 442] = 8'h08; ram[ 443] = 8'h10;
        ram[ 444] = 8'h20; ram[ 445] = 8'h20; ram[ 446] = 8'h20; ram[ 447] = 8'h00;
        ram[ 448] = 8'h38; ram[ 449] = 8'h44; ram[ 450] = 8'h44; ram[ 451] = 8'h38;
        ram[ 452] = 8'h44; ram[ 453] = 8'h44; ram[ 454] = 8'h38; ram[ 455] = 8'h00;
        ram[ 456] = 8'h38; ram[ 457] = 8'h44; ram[ 458] = 8'h44; ram[ 459] = 8'h3C;
        ram[ 460] = 8'h04; ram[ 461] = 8'h08; ram[ 462] = 8'h70; ram[ 463] = 8'h00;
        ram[ 464] = 8'h00; ram[ 465] = 8'h00; ram[ 466] = 8'h10; ram[ 467] = 8'h00;
        ram[ 468] = 8'h10; ram[ 469] = 8'h00; ram[ 470] = 8'h00; ram[ 471] = 8'h00;
        ram[ 472] = 8'h00; ram[ 473] = 8'h00; ram[ 474] = 8'h10; ram[ 475] = 8'h00;
        ram[ 476] = 8'h10; ram[ 477] = 8'h10; ram[ 478] = 8'h20; ram[ 479] = 8'h00;
        ram[ 480] = 8'h08; ram[ 481] = 8'h10; ram[ 482] = 8'h20; ram[ 483] = 8'h40;
        ram[ 484] = 8'h20; ram[ 485] = 8'h10; ram[ 486] = 8'h08; ram[ 487] = 8'h00;
        ram[ 488] = 8'h00; ram[ 489] = 8'h00; ram[ 490] = 8'h7C; ram[ 491] = 8'h00;
        ram[ 492] = 8'h7C; ram[ 493] = 8'h00; ram[ 494] = 8'h00; ram[ 495] = 8'h00;
        ram[ 496] = 8'h20; ram[ 497] = 8'h10; ram[ 498] = 8'h08; ram[ 499] = 8'h04;
        ram[ 500] = 8'h08; ram[ 501] = 8'h10; ram[ 502] = 8'h20; ram[ 503] = 8'h00;
        ram[ 504] = 8'h38; ram[ 505] = 8'h44; ram[ 506] = 8'h08; ram[ 507] = 8'h10;
        ram[ 508] = 8'h10; ram[ 509] = 8'h00; ram[ 510] = 8'h10; ram[ 511] = 8'h00;
        ram[ 512] = 8'h38; ram[ 513] = 8'h44; ram[ 514] = 8'h54; ram[ 515] = 8'h5C;
        ram[ 516] = 8'h58; ram[ 517] = 8'h40; ram[ 518] = 8'h3C; ram[ 519] = 8'h00;
        ram[ 520] = 8'h10; ram[ 521] = 8'h28; ram[ 522] = 8'h44; ram[ 523] = 8'h44;
        ram[ 524] = 8'h7C; ram[ 525] = 8'h44; ram[ 526] = 8'h44; ram[ 527] = 8'h00;
        ram[ 528] = 8'h78; ram[ 529] = 8'h44; ram[ 530] = 8'h44; ram[ 531] = 8'h78;
        ram[ 532] = 8'h44; ram[ 533] = 8'h44; ram[ 534] = 8'h78; ram[ 535] = 8'h00;
        ram[ 536] = 8'h38; ram[ 537] = 8'h44; ram[ 538] = 8'h40; ram[ 539] = 8'h40;
        ram[ 540] = 8'h40; ram[ 541] = 8'h44; ram[ 542] = 8'h38; ram[ 543] = 8'h00;
        ram[ 544] = 8'h78; ram[ 545] = 8'h44; ram[ 546] = 8'h44; ram[ 547] = 8'h44;
        ram[ 548] = 8'h44; ram[ 549] = 8'h44; ram[ 550] = 8'h78; ram[ 551] = 8'h00;
        ram[ 552] = 8'h7C; ram[ 553] = 8'h40; ram[ 554] = 8'h40; ram[ 555] = 8'h78;
        ram[ 556] = 8'h40; ram[ 557] = 8'h40; ram[ 558] = 8'h7C; ram[ 559] = 8'h00;
        ram[ 560] = 8'h7C; ram[ 561] = 8'h40; ram[ 562] = 8'h40; ram[ 563] = 8'h78;
        ram[ 564] = 8'h40; ram[ 565] = 8'h40; ram[ 566] = 8'h40; ram[ 567] = 8'h00;
        ram[ 568] = 8'h3C; ram[ 569] = 8'h40; ram[ 570] = 8'h40; ram[ 571] = 8'h40;
        ram[ 572] = 8'h4C; ram[ 573] = 8'h44; ram[ 574] = 8'h3C; ram[ 575] = 8'h00;
        ram[ 576] = 8'h44; ram[ 577] = 8'h44; ram[ 578] = 8'h44; ram[ 579] = 8'h7C;
        ram[ 580] = 8'h44; ram[ 581] = 8'h44; ram[ 582] = 8'h44; ram[ 583] = 8'h00;
        ram[ 584] = 8'h38; ram[ 585] = 8'h10; ram[ 586] = 8'h10; ram[ 587] = 8'h10;
        ram[ 588] = 8'h10; ram[ 589] = 8'h10; ram[ 590] = 8'h38; ram[ 591] = 8'h00;
        ram[ 592] = 8'h04; ram[ 593] = 8'h04; ram[ 594] = 8'h04; ram[ 595] = 8'h04;
        ram[ 596] = 8'h04; ram[ 597] = 8'h44; ram[ 598] = 8'h38; ram[ 599] = 8'h00;
        ram[ 600] = 8'h44; ram[ 601] = 8'h48; ram[ 602] = 8'h50; ram[ 603] = 8'h60;
        ram[ 604] = 8'h50; ram[ 605] = 8'h48; ram[ 606] = 8'h44; ram[ 607] = 8'h00;
        ram[ 608] = 8'h40; ram[ 609] = 8'h40; ram[ 610] = 8'h40; ram[ 611] = 8'h40;
        ram[ 612] = 8'h40; ram[ 613] = 8'h40; ram[ 614] = 8'h7C; ram[ 615] = 8'h00;
        ram[ 616] = 8'h44; ram[ 617] = 8'h6C; ram[ 618] = 8'h54; ram[ 619] = 8'h54;
        ram[ 620] = 8'h44; ram[ 621] = 8'h44; ram[ 622] = 8'h44; ram[ 623] = 8'h00;
        ram[ 624] = 8'h44; ram[ 625] = 8'h44; ram[ 626] = 8'h64; ram[ 627] = 8'h54;
        ram[ 628] = 8'h4C; ram[ 629] = 8'h44; ram[ 630] = 8'h44; ram[ 631] = 8'h00;
        ram[ 632] = 8'h38; ram[ 633] = 8'h44; ram[ 634] = 8'h44; ram[ 635] = 8'h44;
        ram[ 636] = 8'h44; ram[ 637] = 8'h44; ram[ 638] = 8'h38; ram[ 639] = 8'h00;
        ram[ 640] = 8'h78; ram[ 641] = 8'h44; ram[ 642] = 8'h44; ram[ 643] = 8'h78;
        ram[ 644] = 8'h40; ram[ 645] = 8'h40; ram[ 646] = 8'h40; ram[ 647] = 8'h00;
        ram[ 648] = 8'h38; ram[ 649] = 8'h44; ram[ 650] = 8'h44; ram[ 651] = 8'h44;
        ram[ 652] = 8'h54; ram[ 653] = 8'h48; ram[ 654] = 8'h34; ram[ 655] = 8'h00;
        ram[ 656] = 8'h78; ram[ 657] = 8'h44; ram[ 658] = 8'h44; ram[ 659] = 8'h78;
        ram[ 660] = 8'h50; ram[ 661] = 8'h48; ram[ 662] = 8'h44; ram[ 663] = 8'h00;
        ram[ 664] = 8'h38; ram[ 665] = 8'h44; ram[ 666] = 8'h40; ram[ 667] = 8'h38;
        ram[ 668] = 8'h04; ram[ 669] = 8'h44; ram[ 670] = 8'h38; ram[ 671] = 8'h00;
        ram[ 672] = 8'h7C; ram[ 673] = 8'h10; ram[ 674] = 8'h10; ram[ 675] = 8'h10;
        ram[ 676] = 8'h10; ram[ 677] = 8'h10; ram[ 678] = 8'h10; ram[ 679] = 8'h00;
        ram[ 680] = 8'h44; ram[ 681] = 8'h44; ram[ 682] = 8'h44; ram[ 683] = 8'h44;
        ram[ 684] = 8'h44; ram[ 685] = 8'h44; ram[ 686] = 8'h38; ram[ 687] = 8'h00;
        ram[ 688] = 8'h44; ram[ 689] = 8'h44; ram[ 690] = 8'h44; ram[ 691] = 8'h44;
        ram[ 692] = 8'h44; ram[ 693] = 8'h28; ram[ 694] = 8'h10; ram[ 695] = 8'h00;
        ram[ 696] = 8'h44; ram[ 697] = 8'h44; ram[ 698] = 8'h44; ram[ 699] = 8'h54;
        ram[ 700] = 8'h54; ram[ 701] = 8'h6C; ram[ 702] = 8'h44; ram[ 703] = 8'h00;
        ram[ 704] = 8'h44; ram[ 705] = 8'h44; ram[ 706] = 8'h28; ram[ 707] = 8'h10;
        ram[ 708] = 8'h28; ram[ 709] = 8'h44; ram[ 710] = 8'h44; ram[ 711] = 8'h00;
        ram[ 712] = 8'h44; ram[ 713] = 8'h44; ram[ 714] = 8'h28; ram[ 715] = 8'h10;
        ram[ 716] = 8'h10; ram[ 717] = 8'h10; ram[ 718] = 8'h10; ram[ 719] = 8'h00;
        ram[ 720] = 8'h7C; ram[ 721] = 8'h04; ram[ 722] = 8'h08; ram[ 723] = 8'h10;
        ram[ 724] = 8'h20; ram[ 725] = 8'h40; ram[ 726] = 8'h7C; ram[ 727] = 8'h00;
        ram[ 728] = 8'h7C; ram[ 729] = 8'h60; ram[ 730] = 8'h60; ram[ 731] = 8'h60;
        ram[ 732] = 8'h60; ram[ 733] = 8'h60; ram[ 734] = 8'h7C; ram[ 735] = 8'h00;
        ram[ 736] = 8'h00; ram[ 737] = 8'h40; ram[ 738] = 8'h20; ram[ 739] = 8'h10;
        ram[ 740] = 8'h08; ram[ 741] = 8'h04; ram[ 742] = 8'h00; ram[ 743] = 8'h00;
        ram[ 744] = 8'h7C; ram[ 745] = 8'h0C; ram[ 746] = 8'h0C; ram[ 747] = 8'h0C;
        ram[ 748] = 8'h0C; ram[ 749] = 8'h0C; ram[ 750] = 8'h7C; ram[ 751] = 8'h00;
        ram[ 752] = 8'h00; ram[ 753] = 8'h00; ram[ 754] = 8'h10; ram[ 755] = 8'h28;
        ram[ 756] = 8'h44; ram[ 757] = 8'h00; ram[ 758] = 8'h00; ram[ 759] = 8'h00;
        ram[ 760] = 8'h00; ram[ 761] = 8'h00; ram[ 762] = 8'h00; ram[ 763] = 8'h00;
        ram[ 764] = 8'h00; ram[ 765] = 8'h00; ram[ 766] = 8'h7C; ram[ 767] = 8'h00;
        ram[ 768] = 8'h20; ram[ 769] = 8'h20; ram[ 770] = 8'h10; ram[ 771] = 8'h00;
        ram[ 772] = 8'h00; ram[ 773] = 8'h00; ram[ 774] = 8'h00; ram[ 775] = 8'h00;
        ram[ 776] = 8'h00; ram[ 777] = 8'h00; ram[ 778] = 8'h34; ram[ 779] = 8'h4C;
        ram[ 780] = 8'h44; ram[ 781] = 8'h4C; ram[ 782] = 8'h34; ram[ 783] = 8'h00;
        ram[ 784] = 8'h40; ram[ 785] = 8'h40; ram[ 786] = 8'h58; ram[ 787] = 8'h64;
        ram[ 788] = 8'h44; ram[ 789] = 8'h64; ram[ 790] = 8'h58; ram[ 791] = 8'h00;
        ram[ 792] = 8'h00; ram[ 793] = 8'h00; ram[ 794] = 8'h1C; ram[ 795] = 8'h20;
        ram[ 796] = 8'h20; ram[ 797] = 8'h20; ram[ 798] = 8'h1C; ram[ 799] = 8'h00;
        ram[ 800] = 8'h04; ram[ 801] = 8'h04; ram[ 802] = 8'h34; ram[ 803] = 8'h4C;
        ram[ 804] = 8'h44; ram[ 805] = 8'h4C; ram[ 806] = 8'h34; ram[ 807] = 8'h00;
        ram[ 808] = 8'h00; ram[ 809] = 8'h00; ram[ 810] = 8'h38; ram[ 811] = 8'h44;
        ram[ 812] = 8'h7C; ram[ 813] = 8'h40; ram[ 814] = 8'h38; ram[ 815] = 8'h00;
        ram[ 816] = 8'h08; ram[ 817] = 8'h10; ram[ 818] = 8'h10; ram[ 819] = 8'h38;
        ram[ 820] = 8'h10; ram[ 821] = 8'h10; ram[ 822] = 8'h10; ram[ 823] = 8'h00;
        ram[ 824] = 8'h00; ram[ 825] = 8'h00; ram[ 826] = 8'h34; ram[ 827] = 8'h4C;
        ram[ 828] = 8'h44; ram[ 829] = 8'h3C; ram[ 830] = 8'h04; ram[ 831] = 8'h38;
        ram[ 832] = 8'h40; ram[ 833] = 8'h40; ram[ 834] = 8'h78; ram[ 835] = 8'h44;
        ram[ 836] = 8'h44; ram[ 837] = 8'h44; ram[ 838] = 8'h44; ram[ 839] = 8'h00;
        ram[ 840] = 8'h10; ram[ 841] = 8'h00; ram[ 842] = 8'h30; ram[ 843] = 8'h10;
        ram[ 844] = 8'h10; ram[ 845] = 8'h10; ram[ 846] = 8'h38; ram[ 847] = 8'h00;
        ram[ 848] = 8'h08; ram[ 849] = 8'h00; ram[ 850] = 8'h08; ram[ 851] = 8'h08;
        ram[ 852] = 8'h08; ram[ 853] = 8'h08; ram[ 854] = 8'h08; ram[ 855] = 8'h30;
        ram[ 856] = 8'h40; ram[ 857] = 8'h40; ram[ 858] = 8'h48; ram[ 859] = 8'h50;
        ram[ 860] = 8'h70; ram[ 861] = 8'h48; ram[ 862] = 8'h44; ram[ 863] = 8'h00;
        ram[ 864] = 8'h30; ram[ 865] = 8'h10; ram[ 866] = 8'h10; ram[ 867] = 8'h10;
        ram[ 868] = 8'h10; ram[ 869] = 8'h10; ram[ 870] = 8'h38; ram[ 871] = 8'h00;
        ram[ 872] = 8'h00; ram[ 873] = 8'h00; ram[ 874] = 8'h6C; ram[ 875] = 8'h52;
        ram[ 876] = 8'h52; ram[ 877] = 8'h52; ram[ 878] = 8'h52; ram[ 879] = 8'h00;
        ram[ 880] = 8'h00; ram[ 881] = 8'h00; ram[ 882] = 8'h78; ram[ 883] = 8'h44;
        ram[ 884] = 8'h44; ram[ 885] = 8'h44; ram[ 886] = 8'h44; ram[ 887] = 8'h00;
        ram[ 888] = 8'h00; ram[ 889] = 8'h00; ram[ 890] = 8'h38; ram[ 891] = 8'h44;
        ram[ 892] = 8'h44; ram[ 893] = 8'h44; ram[ 894] = 8'h38; ram[ 895] = 8'h00;
        ram[ 896] = 8'h00; ram[ 897] = 8'h00; ram[ 898] = 8'h58; ram[ 899] = 8'h64;
        ram[ 900] = 8'h44; ram[ 901] = 8'h64; ram[ 902] = 8'h58; ram[ 903] = 8'h40;
        ram[ 904] = 8'h00; ram[ 905] = 8'h00; ram[ 906] = 8'h34; ram[ 907] = 8'h4C;
        ram[ 908] = 8'h44; ram[ 909] = 8'h4C; ram[ 910] = 8'h34; ram[ 911] = 8'h06;
        ram[ 912] = 8'h00; ram[ 913] = 8'h00; ram[ 914] = 8'h58; ram[ 915] = 8'h60;
        ram[ 916] = 8'h40; ram[ 917] = 8'h40; ram[ 918] = 8'h40; ram[ 919] = 8'h00;
        ram[ 920] = 8'h00; ram[ 921] = 8'h00; ram[ 922] = 8'h3C; ram[ 923] = 8'h40;
        ram[ 924] = 8'h38; ram[ 925] = 8'h04; ram[ 926] = 8'h78; ram[ 927] = 8'h00;
        ram[ 928] = 8'h10; ram[ 929] = 8'h10; ram[ 930] = 8'h7C; ram[ 931] = 8'h10;
        ram[ 932] = 8'h10; ram[ 933] = 8'h10; ram[ 934] = 8'h10; ram[ 935] = 8'h00;
        ram[ 936] = 8'h00; ram[ 937] = 8'h00; ram[ 938] = 8'h44; ram[ 939] = 8'h44;
        ram[ 940] = 8'h44; ram[ 941] = 8'h44; ram[ 942] = 8'h3C; ram[ 943] = 8'h00;
        ram[ 944] = 8'h00; ram[ 945] = 8'h00; ram[ 946] = 8'h44; ram[ 947] = 8'h44;
        ram[ 948] = 8'h28; ram[ 949] = 8'h28; ram[ 950] = 8'h10; ram[ 951] = 8'h00;
        ram[ 952] = 8'h00; ram[ 953] = 8'h00; ram[ 954] = 8'h52; ram[ 955] = 8'h52;
        ram[ 956] = 8'h52; ram[ 957] = 8'h52; ram[ 958] = 8'h2C; ram[ 959] = 8'h00;
        ram[ 960] = 8'h00; ram[ 961] = 8'h00; ram[ 962] = 8'h44; ram[ 963] = 8'h28;
        ram[ 964] = 8'h10; ram[ 965] = 8'h28; ram[ 966] = 8'h44; ram[ 967] = 8'h00;
        ram[ 968] = 8'h00; ram[ 969] = 8'h00; ram[ 970] = 8'h24; ram[ 971] = 8'h24;
        ram[ 972] = 8'h24; ram[ 973] = 8'h3C; ram[ 974] = 8'h04; ram[ 975] = 8'h38;
        ram[ 976] = 8'h00; ram[ 977] = 8'h00; ram[ 978] = 8'h7C; ram[ 979] = 8'h08;
        ram[ 980] = 8'h10; ram[ 981] = 8'h20; ram[ 982] = 8'h7C; ram[ 983] = 8'h00;
        ram[ 984] = 8'h0C; ram[ 985] = 8'h10; ram[ 986] = 8'h10; ram[ 987] = 8'h20;
        ram[ 988] = 8'h10; ram[ 989] = 8'h10; ram[ 990] = 8'h0C; ram[ 991] = 8'h00;
        ram[ 992] = 8'h10; ram[ 993] = 8'h10; ram[ 994] = 8'h10; ram[ 995] = 8'h00;
        ram[ 996] = 8'h10; ram[ 997] = 8'h10; ram[ 998] = 8'h10; ram[ 999] = 8'h00;
        ram[1000] = 8'h60; ram[1001] = 8'h10; ram[1002] = 8'h10; ram[1003] = 8'h08;
        ram[1004] = 8'h10; ram[1005] = 8'h10; ram[1006] = 8'h60; ram[1007] = 8'h00;
        ram[1008] = 8'h00; ram[1009] = 8'h00; ram[1010] = 8'h04; ram[1011] = 8'h38;
        ram[1012] = 8'h40; ram[1013] = 8'h00; ram[1014] = 8'h00; ram[1015] = 8'h00;
        ram[1016] = 8'hFF; ram[1017] = 8'hFF; ram[1018] = 8'hFF; ram[1019] = 8'hFF;
        ram[1020] = 8'hFF; ram[1021] = 8'hFF; ram[1022] = 8'hFF; ram[1023] = 8'hFF;
        ram[1024] = 8'h00; ram[1025] = 8'hFF; ram[1026] = 8'hFF; ram[1027] = 8'hFF;
        ram[1028] = 8'hFF; ram[1029] = 8'hFF; ram[1030] = 8'hFF; ram[1031] = 8'hFF;
        ram[1032] = 8'h80; ram[1033] = 8'h80; ram[1034] = 8'h80; ram[1035] = 8'h80;
        ram[1036] = 8'h80; ram[1037] = 8'h80; ram[1038] = 8'h80; ram[1039] = 8'h80;
        ram[1040] = 8'h00; ram[1041] = 8'h1C; ram[1042] = 8'h3C; ram[1043] = 8'h00;
        ram[1044] = 8'h1C; ram[1045] = 8'h1E; ram[1046] = 8'h3E; ram[1047] = 8'hFE;
        ram[1048] = 8'h3E; ram[1049] = 8'h7C; ram[1050] = 8'hD8; ram[1051] = 8'h78;
        ram[1052] = 8'h38; ram[1053] = 8'h18; ram[1054] = 8'h1C; ram[1055] = 8'h1C;
        ram[1056] = 8'h00; ram[1057] = 8'h00; ram[1058] = 8'h00; ram[1059] = 8'h00;
        ram[1060] = 8'hAA; ram[1061] = 8'h55; ram[1062] = 8'hAA; ram[1063] = 8'h55;
        ram[1064] = 8'hA0; ram[1065] = 8'h50; ram[1066] = 8'hA0; ram[1067] = 8'h50;
        ram[1068] = 8'hA0; ram[1069] = 8'h50; ram[1070] = 8'hA0; ram[1071] = 8'h50;
        ram[1072] = 8'hAA; ram[1073] = 8'h55; ram[1074] = 8'hAA; ram[1075] = 8'h55;
        ram[1076] = 8'hAA; ram[1077] = 8'h55; ram[1078] = 8'hAA; ram[1079] = 8'h55;
        ram[1080] = 8'h00; ram[1081] = 8'h18; ram[1082] = 8'h3C; ram[1083] = 8'h7E;
        ram[1084] = 8'h7E; ram[1085] = 8'h3C; ram[1086] = 8'h18; ram[1087] = 8'h00;
        ram[1088] = 8'h00; ram[1089] = 8'h00; ram[1090] = 8'h00; ram[1091] = 8'h00;
        ram[1092] = 8'h00; ram[1093] = 8'h00; ram[1094] = 8'hFF; ram[1095] = 8'hFF;
        ram[1096] = 8'h00; ram[1097] = 8'h00; ram[1098] = 8'hFF; ram[1099] = 8'hFF;
        ram[1100] = 8'hFF; ram[1101] = 8'hFF; ram[1102] = 8'hFF; ram[1103] = 8'hFF;
        ram[1104] = 8'h18; ram[1105] = 8'h18; ram[1106] = 8'h3C; ram[1107] = 8'h7E;
        ram[1108] = 8'hFF; ram[1109] = 8'hDB; ram[1110] = 8'h18; ram[1111] = 8'h3C;
        ram[1112] = 8'h3C; ram[1113] = 8'h18; ram[1114] = 8'hDB; ram[1115] = 8'hFF;
        ram[1116] = 8'h7E; ram[1117] = 8'h3C; ram[1118] = 8'h18; ram[1119] = 8'h18;
        ram[1120] = 8'h00; ram[1121] = 8'h1C; ram[1122] = 8'h3C; ram[1123] = 8'h00;
        ram[1124] = 8'h9C; ram[1125] = 8'h9E; ram[1126] = 8'hFB; ram[1127] = 8'h3B;
        ram[1128] = 8'h3E; ram[1129] = 8'hFC; ram[1130] = 8'hF8; ram[1131] = 8'hDC;
        ram[1132] = 8'hCF; ram[1133] = 8'hC3; ram[1134] = 8'h01; ram[1135] = 8'h00;
        ram[1136] = 8'hC0; ram[1137] = 8'hF0; ram[1138] = 8'hFC; ram[1139] = 8'hFF;
        ram[1140] = 8'hFF; ram[1141] = 8'hFC; ram[1142] = 8'hF0; ram[1143] = 8'hC0;
        ram[1144] = 8'h18; ram[1145] = 8'h18; ram[1146] = 8'h3C; ram[1147] = 8'h3C;
        ram[1148] = 8'h7E; ram[1149] = 8'h7E; ram[1150] = 8'hFF; ram[1151] = 8'hFF;
        ram[1152] = 8'h00; ram[1153] = 8'h00; ram[1154] = 8'h00; ram[1155] = 8'h00;
        ram[1156] = 8'h00; ram[1157] = 8'h00; ram[1158] = 8'h00; ram[1159] = 8'hFF;
        ram[1160] = 8'hFE; ram[1161] = 8'hFE; ram[1162] = 8'hFE; ram[1163] = 8'hFE;
        ram[1164] = 8'hFE; ram[1165] = 8'hFE; ram[1166] = 8'hFE; ram[1167] = 8'hFE;
        ram[1168] = 8'h3C; ram[1169] = 8'h52; ram[1170] = 8'h3C; ram[1171] = 8'h80;
        ram[1172] = 8'hBC; ram[1173] = 8'hFF; ram[1174] = 8'h3D; ram[1175] = 8'h3D;
        ram[1176] = 8'h3C; ram[1177] = 8'h4A; ram[1178] = 8'h3C; ram[1179] = 8'h01;
        ram[1180] = 8'h3D; ram[1181] = 8'hFF; ram[1182] = 8'hBC; ram[1183] = 8'hBC;
        ram[1184] = 8'hAA; ram[1185] = 8'h55; ram[1186] = 8'hAA; ram[1187] = 8'h55;
        ram[1188] = 8'h00; ram[1189] = 8'h00; ram[1190] = 8'h00; ram[1191] = 8'h00;
        ram[1192] = 8'h0A; ram[1193] = 8'h05; ram[1194] = 8'h0A; ram[1195] = 8'h05;
        ram[1196] = 8'h0A; ram[1197] = 8'h05; ram[1198] = 8'h0A; ram[1199] = 8'h05;
        ram[1200] = 8'h3C; ram[1201] = 8'h7E; ram[1202] = 8'hFF; ram[1203] = 8'hFF;
        ram[1204] = 8'hFF; ram[1205] = 8'hFF; ram[1206] = 8'h7E; ram[1207] = 8'h3C;
        ram[1208] = 8'hC0; ram[1209] = 8'hC0; ram[1210] = 8'hC0; ram[1211] = 8'hC0;
        ram[1212] = 8'hC0; ram[1213] = 8'hC0; ram[1214] = 8'hC0; ram[1215] = 8'hC0;
        ram[1216] = 8'hE0; ram[1217] = 8'hE0; ram[1218] = 8'hE0; ram[1219] = 8'hE0;
        ram[1220] = 8'hE0; ram[1221] = 8'hE0; ram[1222] = 8'hE0; ram[1223] = 8'hE0;
        ram[1224] = 8'hF8; ram[1225] = 8'hF8; ram[1226] = 8'hF8; ram[1227] = 8'hF8;
        ram[1228] = 8'hF8; ram[1229] = 8'hF8; ram[1230] = 8'hF8; ram[1231] = 8'hF8;
        ram[1232] = 8'h30; ram[1233] = 8'h38; ram[1234] = 8'h9C; ram[1235] = 8'hFF;
        ram[1236] = 8'hFF; ram[1237] = 8'h9C; ram[1238] = 8'h38; ram[1239] = 8'h30;
        ram[1240] = 8'h0C; ram[1241] = 8'h1C; ram[1242] = 8'h39; ram[1243] = 8'hFF;
        ram[1244] = 8'hFF; ram[1245] = 8'h39; ram[1246] = 8'h1C; ram[1247] = 8'h0C;
        ram[1248] = 8'h00; ram[1249] = 8'h66; ram[1250] = 8'h7E; ram[1251] = 8'h42;
        ram[1252] = 8'hC3; ram[1253] = 8'hFF; ram[1254] = 8'h18; ram[1255] = 8'h00;
        ram[1256] = 8'h00; ram[1257] = 8'h18; ram[1258] = 8'hFF; ram[1259] = 8'hC3;
        ram[1260] = 8'h42; ram[1261] = 8'h7E; ram[1262] = 8'h66; ram[1263] = 8'h00;
        ram[1264] = 8'h03; ram[1265] = 8'h0F; ram[1266] = 8'h3F; ram[1267] = 8'hFF;
        ram[1268] = 8'hFF; ram[1269] = 8'h3F; ram[1270] = 8'h0F; ram[1271] = 8'h03;
        ram[1272] = 8'hFF; ram[1273] = 8'hFF; ram[1274] = 8'h7E; ram[1275] = 8'h7E;
        ram[1276] = 8'h3C; ram[1277] = 8'h3C; ram[1278] = 8'h18; ram[1279] = 8'h18;
        ram[1280] = 8'h00; ram[1281] = 8'h00; ram[1282] = 8'h00; ram[1283] = 8'h00;
        ram[1284] = 8'h00; ram[1285] = 8'h00; ram[1286] = 8'h00; ram[1287] = 8'h00;
        ram[1288] = 8'hF0; ram[1289] = 8'hF0; ram[1290] = 8'hF0; ram[1291] = 8'h00;
        ram[1292] = 8'h00; ram[1293] = 8'h00; ram[1294] = 8'h00; ram[1295] = 8'h00;
        ram[1296] = 8'h0F; ram[1297] = 8'h0F; ram[1298] = 8'h0F; ram[1299] = 8'h00;
        ram[1300] = 8'h00; ram[1301] = 8'h00; ram[1302] = 8'h00; ram[1303] = 8'h00;
        ram[1304] = 8'hFF; ram[1305] = 8'hFF; ram[1306] = 8'hFF; ram[1307] = 8'h00;
        ram[1308] = 8'h00; ram[1309] = 8'h00; ram[1310] = 8'h00; ram[1311] = 8'h00;
        ram[1312] = 8'h00; ram[1313] = 8'h00; ram[1314] = 8'h00; ram[1315] = 8'hF0;
        ram[1316] = 8'hF0; ram[1317] = 8'h00; ram[1318] = 8'h00; ram[1319] = 8'h00;
        ram[1320] = 8'hF0; ram[1321] = 8'hF0; ram[1322] = 8'hF0; ram[1323] = 8'hF0;
        ram[1324] = 8'hF0; ram[1325] = 8'h00; ram[1326] = 8'h00; ram[1327] = 8'h00;
        ram[1328] = 8'h0F; ram[1329] = 8'h0F; ram[1330] = 8'h0F; ram[1331] = 8'hF0;
        ram[1332] = 8'hF0; ram[1333] = 8'h00; ram[1334] = 8'h00; ram[1335] = 8'h00;
        ram[1336] = 8'hFF; ram[1337] = 8'hFF; ram[1338] = 8'hFF; ram[1339] = 8'hF0;
        ram[1340] = 8'hF0; ram[1341] = 8'h00; ram[1342] = 8'h00; ram[1343] = 8'h00;
        ram[1344] = 8'h00; ram[1345] = 8'h00; ram[1346] = 8'h00; ram[1347] = 8'h0F;
        ram[1348] = 8'h0F; ram[1349] = 8'h00; ram[1350] = 8'h00; ram[1351] = 8'h00;
        ram[1352] = 8'hF0; ram[1353] = 8'hF0; ram[1354] = 8'hF0; ram[1355] = 8'h0F;
        ram[1356] = 8'h0F; ram[1357] = 8'h00; ram[1358] = 8'h00; ram[1359] = 8'h00;
        ram[1360] = 8'h0F; ram[1361] = 8'h0F; ram[1362] = 8'h0F; ram[1363] = 8'h0F;
        ram[1364] = 8'h0F; ram[1365] = 8'h00; ram[1366] = 8'h00; ram[1367] = 8'h00;
        ram[1368] = 8'hFF; ram[1369] = 8'hFF; ram[1370] = 8'hFF; ram[1371] = 8'h0F;
        ram[1372] = 8'h0F; ram[1373] = 8'h00; ram[1374] = 8'h00; ram[1375] = 8'h00;
        ram[1376] = 8'h00; ram[1377] = 8'h00; ram[1378] = 8'h00; ram[1379] = 8'hFF;
        ram[1380] = 8'hFF; ram[1381] = 8'h00; ram[1382] = 8'h00; ram[1383] = 8'h00;
        ram[1384] = 8'hF0; ram[1385] = 8'hF0; ram[1386] = 8'hF0; ram[1387] = 8'hFF;
        ram[1388] = 8'hFF; ram[1389] = 8'h00; ram[1390] = 8'h00; ram[1391] = 8'h00;
        ram[1392] = 8'h0F; ram[1393] = 8'h0F; ram[1394] = 8'h0F; ram[1395] = 8'hFF;
        ram[1396] = 8'hFF; ram[1397] = 8'h00; ram[1398] = 8'h00; ram[1399] = 8'h00;
        ram[1400] = 8'hFF; ram[1401] = 8'hFF; ram[1402] = 8'hFF; ram[1403] = 8'hFF;
        ram[1404] = 8'hFF; ram[1405] = 8'h00; ram[1406] = 8'h00; ram[1407] = 8'h00;
        ram[1408] = 8'h00; ram[1409] = 8'h00; ram[1410] = 8'h00; ram[1411] = 8'h00;
        ram[1412] = 8'h00; ram[1413] = 8'hF0; ram[1414] = 8'hF0; ram[1415] = 8'hF0;
        ram[1416] = 8'hF0; ram[1417] = 8'hF0; ram[1418] = 8'hF0; ram[1419] = 8'h00;
        ram[1420] = 8'h00; ram[1421] = 8'hF0; ram[1422] = 8'hF0; ram[1423] = 8'hF0;
        ram[1424] = 8'h0F; ram[1425] = 8'h0F; ram[1426] = 8'h0F; ram[1427] = 8'h00;
        ram[1428] = 8'h00; ram[1429] = 8'hF0; ram[1430] = 8'hF0; ram[1431] = 8'hF0;
        ram[1432] = 8'hFF; ram[1433] = 8'hFF; ram[1434] = 8'hFF; ram[1435] = 8'h00;
        ram[1436] = 8'h00; ram[1437] = 8'hF0; ram[1438] = 8'hF0; ram[1439] = 8'hF0;
        ram[1440] = 8'h00; ram[1441] = 8'h00; ram[1442] = 8'h00; ram[1443] = 8'hF0;
        ram[1444] = 8'hF0; ram[1445] = 8'hF0; ram[1446] = 8'hF0; ram[1447] = 8'hF0;
        ram[1448] = 8'hF0; ram[1449] = 8'hF0; ram[1450] = 8'hF0; ram[1451] = 8'hF0;
        ram[1452] = 8'hF0; ram[1453] = 8'hF0; ram[1454] = 8'hF0; ram[1455] = 8'hF0;
        ram[1456] = 8'h0F; ram[1457] = 8'h0F; ram[1458] = 8'h0F; ram[1459] = 8'hF0;
        ram[1460] = 8'hF0; ram[1461] = 8'hF0; ram[1462] = 8'hF0; ram[1463] = 8'hF0;
        ram[1464] = 8'hFF; ram[1465] = 8'hFF; ram[1466] = 8'hFF; ram[1467] = 8'hF0;
        ram[1468] = 8'hF0; ram[1469] = 8'hF0; ram[1470] = 8'hF0; ram[1471] = 8'hF0;
        ram[1472] = 8'h00; ram[1473] = 8'h00; ram[1474] = 8'h00; ram[1475] = 8'h0F;
        ram[1476] = 8'h0F; ram[1477] = 8'hF0; ram[1478] = 8'hF0; ram[1479] = 8'hF0;
        ram[1480] = 8'hF0; ram[1481] = 8'hF0; ram[1482] = 8'hF0; ram[1483] = 8'h0F;
        ram[1484] = 8'h0F; ram[1485] = 8'hF0; ram[1486] = 8'hF0; ram[1487] = 8'hF0;
        ram[1488] = 8'h0F; ram[1489] = 8'h0F; ram[1490] = 8'h0F; ram[1491] = 8'h0F;
        ram[1492] = 8'h0F; ram[1493] = 8'hF0; ram[1494] = 8'hF0; ram[1495] = 8'hF0;
        ram[1496] = 8'hFF; ram[1497] = 8'hFF; ram[1498] = 8'hFF; ram[1499] = 8'h0F;
        ram[1500] = 8'h0F; ram[1501] = 8'hF0; ram[1502] = 8'hF0; ram[1503] = 8'hF0;
        ram[1504] = 8'h00; ram[1505] = 8'h00; ram[1506] = 8'h00; ram[1507] = 8'hFF;
        ram[1508] = 8'hFF; ram[1509] = 8'hF0; ram[1510] = 8'hF0; ram[1511] = 8'hF0;
        ram[1512] = 8'hF0; ram[1513] = 8'hF0; ram[1514] = 8'hF0; ram[1515] = 8'hFF;
        ram[1516] = 8'hFF; ram[1517] = 8'hF0; ram[1518] = 8'hF0; ram[1519] = 8'hF0;
        ram[1520] = 8'h0F; ram[1521] = 8'h0F; ram[1522] = 8'h0F; ram[1523] = 8'hFF;
        ram[1524] = 8'hFF; ram[1525] = 8'hF0; ram[1526] = 8'hF0; ram[1527] = 8'hF0;
        ram[1528] = 8'hFF; ram[1529] = 8'hFF; ram[1530] = 8'hFF; ram[1531] = 8'hFF;
        ram[1532] = 8'hFF; ram[1533] = 8'hF0; ram[1534] = 8'hF0; ram[1535] = 8'hF0;
        ram[1536] = 8'h01; ram[1537] = 8'h03; ram[1538] = 8'h07; ram[1539] = 8'h0F;
        ram[1540] = 8'h1F; ram[1541] = 8'h3F; ram[1542] = 8'h7F; ram[1543] = 8'hFF;
        ram[1544] = 8'h80; ram[1545] = 8'hC0; ram[1546] = 8'hE0; ram[1547] = 8'hF0;
        ram[1548] = 8'hF8; ram[1549] = 8'hFC; ram[1550] = 8'hFE; ram[1551] = 8'hFF;
        ram[1552] = 8'hFF; ram[1553] = 8'hFF; ram[1554] = 8'h7E; ram[1555] = 8'h3C;
        ram[1556] = 8'h00; ram[1557] = 8'h00; ram[1558] = 8'h00; ram[1559] = 8'h00;
        ram[1560] = 8'hFC; ram[1561] = 8'hFC; ram[1562] = 8'hFC; ram[1563] = 8'hFC;
        ram[1564] = 8'hFC; ram[1565] = 8'hFC; ram[1566] = 8'hFC; ram[1567] = 8'hFC;
        ram[1568] = 8'h00; ram[1569] = 8'h00; ram[1570] = 8'h3C; ram[1571] = 8'h3C;
        ram[1572] = 8'h3C; ram[1573] = 8'h3C; ram[1574] = 8'h00; ram[1575] = 8'h00;
        ram[1576] = 8'h18; ram[1577] = 8'h3C; ram[1578] = 8'h7E; ram[1579] = 8'hFF;
        ram[1580] = 8'hFF; ram[1581] = 8'h7E; ram[1582] = 8'h3C; ram[1583] = 8'h18;
        ram[1584] = 8'h00; ram[1585] = 8'h00; ram[1586] = 8'h00; ram[1587] = 8'h18;
        ram[1588] = 8'h18; ram[1589] = 8'h00; ram[1590] = 8'h00; ram[1591] = 8'h00;
        ram[1592] = 8'h0F; ram[1593] = 8'h0F; ram[1594] = 8'h07; ram[1595] = 8'h03;
        ram[1596] = 8'h00; ram[1597] = 8'h00; ram[1598] = 8'h00; ram[1599] = 8'h00;
        ram[1600] = 8'h18; ram[1601] = 8'h18; ram[1602] = 8'h18; ram[1603] = 8'hFF;
        ram[1604] = 8'hFF; ram[1605] = 8'h18; ram[1606] = 8'h18; ram[1607] = 8'h18;
        ram[1608] = 8'h00; ram[1609] = 8'h00; ram[1610] = 8'h00; ram[1611] = 8'h00;
        ram[1612] = 8'hC0; ram[1613] = 8'hE0; ram[1614] = 8'hF0; ram[1615] = 8'hF0;
        ram[1616] = 8'h01; ram[1617] = 8'h02; ram[1618] = 8'h04; ram[1619] = 8'h08;
        ram[1620] = 8'h10; ram[1621] = 8'h20; ram[1622] = 8'h40; ram[1623] = 8'h80;
        ram[1624] = 8'h03; ram[1625] = 8'h07; ram[1626] = 8'h0F; ram[1627] = 8'h0F;
        ram[1628] = 8'h0F; ram[1629] = 8'h0F; ram[1630] = 8'h07; ram[1631] = 8'h03;
        ram[1632] = 8'h18; ram[1633] = 8'h18; ram[1634] = 8'h18; ram[1635] = 8'hFF;
        ram[1636] = 8'hFF; ram[1637] = 8'h00; ram[1638] = 8'h00; ram[1639] = 8'h00;
        ram[1640] = 8'h18; ram[1641] = 8'h18; ram[1642] = 8'h18; ram[1643] = 8'h1F;
        ram[1644] = 8'h1F; ram[1645] = 8'h18; ram[1646] = 8'h18; ram[1647] = 8'h18;
        ram[1648] = 8'h00; ram[1649] = 8'h00; ram[1650] = 8'h00; ram[1651] = 8'hF8;
        ram[1652] = 8'hF8; ram[1653] = 8'h18; ram[1654] = 8'h18; ram[1655] = 8'h18;
        ram[1656] = 8'h18; ram[1657] = 8'h18; ram[1658] = 8'h18; ram[1659] = 8'h1F;
        ram[1660] = 8'h1F; ram[1661] = 8'h00; ram[1662] = 8'h00; ram[1663] = 8'h00;
        ram[1664] = 8'h09; ram[1665] = 8'h20; ram[1666] = 8'h04; ram[1667] = 8'h80;
        ram[1668] = 8'h11; ram[1669] = 8'h40; ram[1670] = 8'h08; ram[1671] = 8'h02;
        ram[1672] = 8'h52; ram[1673] = 8'h44; ram[1674] = 8'h2D; ram[1675] = 8'hC4;
        ram[1676] = 8'h11; ram[1677] = 8'hB4; ram[1678] = 8'h23; ram[1679] = 8'h4A;
        ram[1680] = 8'h00; ram[1681] = 8'h00; ram[1682] = 8'h00; ram[1683] = 8'h00;
        ram[1684] = 8'h3C; ram[1685] = 8'h7E; ram[1686] = 8'hFF; ram[1687] = 8'hFF;
        ram[1688] = 8'h00; ram[1689] = 8'h10; ram[1690] = 8'h2C; ram[1691] = 8'h3A;
        ram[1692] = 8'h5C; ram[1693] = 8'h34; ram[1694] = 8'h04; ram[1695] = 8'h00;
        ram[1696] = 8'h66; ram[1697] = 8'hFF; ram[1698] = 8'hFF; ram[1699] = 8'hFF;
        ram[1700] = 8'h7E; ram[1701] = 8'h3C; ram[1702] = 8'h18; ram[1703] = 8'h18;
        ram[1704] = 8'h18; ram[1705] = 8'h3C; ram[1706] = 8'h18; ram[1707] = 8'h42;
        ram[1708] = 8'hE7; ram[1709] = 8'h42; ram[1710] = 8'h18; ram[1711] = 8'h3C;
        ram[1712] = 8'h18; ram[1713] = 8'h18; ram[1714] = 8'h18; ram[1715] = 8'h18;
        ram[1716] = 8'h18; ram[1717] = 8'h18; ram[1718] = 8'h18; ram[1719] = 8'h18;
        ram[1720] = 8'h00; ram[1721] = 8'h00; ram[1722] = 8'h00; ram[1723] = 8'h00;
        ram[1724] = 8'h03; ram[1725] = 8'h07; ram[1726] = 8'h0F; ram[1727] = 8'h0F;
        ram[1728] = 8'h81; ram[1729] = 8'h42; ram[1730] = 8'h24; ram[1731] = 8'h18;
        ram[1732] = 8'h18; ram[1733] = 8'h24; ram[1734] = 8'h42; ram[1735] = 8'h81;
        ram[1736] = 8'hF0; ram[1737] = 8'hF0; ram[1738] = 8'hE0; ram[1739] = 8'hC0;
        ram[1740] = 8'h00; ram[1741] = 8'h00; ram[1742] = 8'h00; ram[1743] = 8'h00;
        ram[1744] = 8'h80; ram[1745] = 8'h40; ram[1746] = 8'h20; ram[1747] = 8'h10;
        ram[1748] = 8'h08; ram[1749] = 8'h04; ram[1750] = 8'h02; ram[1751] = 8'h01;
        ram[1752] = 8'hC0; ram[1753] = 8'hE0; ram[1754] = 8'hF0; ram[1755] = 8'hF0;
        ram[1756] = 8'hF0; ram[1757] = 8'hF0; ram[1758] = 8'hE0; ram[1759] = 8'hC0;
        ram[1760] = 8'h00; ram[1761] = 8'h00; ram[1762] = 8'h00; ram[1763] = 8'hFF;
        ram[1764] = 8'hFF; ram[1765] = 8'h18; ram[1766] = 8'h18; ram[1767] = 8'h18;
        ram[1768] = 8'h18; ram[1769] = 8'h18; ram[1770] = 8'h18; ram[1771] = 8'hF8;
        ram[1772] = 8'hF8; ram[1773] = 8'h18; ram[1774] = 8'h18; ram[1775] = 8'h18;
        ram[1776] = 8'h00; ram[1777] = 8'h00; ram[1778] = 8'h00; ram[1779] = 8'h1F;
        ram[1780] = 8'h1F; ram[1781] = 8'h18; ram[1782] = 8'h18; ram[1783] = 8'h18;
        ram[1784] = 8'h18; ram[1785] = 8'h18; ram[1786] = 8'h18; ram[1787] = 8'hF8;
        ram[1788] = 8'hF8; ram[1789] = 8'h00; ram[1790] = 8'h00; ram[1791] = 8'h00;
        ram[1792] = 8'h00; ram[1793] = 8'h00; ram[1794] = 8'h00; ram[1795] = 8'h00;
        ram[1796] = 8'h00; ram[1797] = 8'h0F; ram[1798] = 8'h0F; ram[1799] = 8'h0F;
        ram[1800] = 8'hF0; ram[1801] = 8'hF0; ram[1802] = 8'hF0; ram[1803] = 8'h00;
        ram[1804] = 8'h00; ram[1805] = 8'h0F; ram[1806] = 8'h0F; ram[1807] = 8'h0F;
        ram[1808] = 8'h0F; ram[1809] = 8'h0F; ram[1810] = 8'h0F; ram[1811] = 8'h00;
        ram[1812] = 8'h00; ram[1813] = 8'h0F; ram[1814] = 8'h0F; ram[1815] = 8'h0F;
        ram[1816] = 8'hFF; ram[1817] = 8'hFF; ram[1818] = 8'hFF; ram[1819] = 8'h00;
        ram[1820] = 8'h00; ram[1821] = 8'h0F; ram[1822] = 8'h0F; ram[1823] = 8'h0F;
        ram[1824] = 8'h00; ram[1825] = 8'h00; ram[1826] = 8'h00; ram[1827] = 8'hF0;
        ram[1828] = 8'hF0; ram[1829] = 8'h0F; ram[1830] = 8'h0F; ram[1831] = 8'h0F;
        ram[1832] = 8'hF0; ram[1833] = 8'hF0; ram[1834] = 8'hF0; ram[1835] = 8'hF0;
        ram[1836] = 8'hF0; ram[1837] = 8'h0F; ram[1838] = 8'h0F; ram[1839] = 8'h0F;
        ram[1840] = 8'h0F; ram[1841] = 8'h0F; ram[1842] = 8'h0F; ram[1843] = 8'hF0;
        ram[1844] = 8'hF0; ram[1845] = 8'h0F; ram[1846] = 8'h0F; ram[1847] = 8'h0F;
        ram[1848] = 8'hFF; ram[1849] = 8'hFF; ram[1850] = 8'hFF; ram[1851] = 8'hF0;
        ram[1852] = 8'hF0; ram[1853] = 8'h0F; ram[1854] = 8'h0F; ram[1855] = 8'h0F;
        ram[1856] = 8'h00; ram[1857] = 8'h00; ram[1858] = 8'h00; ram[1859] = 8'h0F;
        ram[1860] = 8'h0F; ram[1861] = 8'h0F; ram[1862] = 8'h0F; ram[1863] = 8'h0F;
        ram[1864] = 8'hF0; ram[1865] = 8'hF0; ram[1866] = 8'hF0; ram[1867] = 8'h0F;
        ram[1868] = 8'h0F; ram[1869] = 8'h0F; ram[1870] = 8'h0F; ram[1871] = 8'h0F;
        ram[1872] = 8'h0F; ram[1873] = 8'h0F; ram[1874] = 8'h0F; ram[1875] = 8'h0F;
        ram[1876] = 8'h0F; ram[1877] = 8'h0F; ram[1878] = 8'h0F; ram[1879] = 8'h0F;
        ram[1880] = 8'hFF; ram[1881] = 8'hFF; ram[1882] = 8'hFF; ram[1883] = 8'h0F;
        ram[1884] = 8'h0F; ram[1885] = 8'h0F; ram[1886] = 8'h0F; ram[1887] = 8'h0F;
        ram[1888] = 8'h00; ram[1889] = 8'h00; ram[1890] = 8'h00; ram[1891] = 8'hFF;
        ram[1892] = 8'hFF; ram[1893] = 8'h0F; ram[1894] = 8'h0F; ram[1895] = 8'h0F;
        ram[1896] = 8'hF0; ram[1897] = 8'hF0; ram[1898] = 8'hF0; ram[1899] = 8'hFF;
        ram[1900] = 8'hFF; ram[1901] = 8'h0F; ram[1902] = 8'h0F; ram[1903] = 8'h0F;
        ram[1904] = 8'h0F; ram[1905] = 8'h0F; ram[1906] = 8'h0F; ram[1907] = 8'hFF;
        ram[1908] = 8'hFF; ram[1909] = 8'h0F; ram[1910] = 8'h0F; ram[1911] = 8'h0F;
        ram[1912] = 8'hFF; ram[1913] = 8'hFF; ram[1914] = 8'hFF; ram[1915] = 8'hFF;
        ram[1916] = 8'hFF; ram[1917] = 8'h0F; ram[1918] = 8'h0F; ram[1919] = 8'h0F;
        ram[1920] = 8'h00; ram[1921] = 8'h00; ram[1922] = 8'h00; ram[1923] = 8'h00;
        ram[1924] = 8'h00; ram[1925] = 8'hFF; ram[1926] = 8'hFF; ram[1927] = 8'hFF;
        ram[1928] = 8'hF0; ram[1929] = 8'hF0; ram[1930] = 8'hF0; ram[1931] = 8'h00;
        ram[1932] = 8'h00; ram[1933] = 8'hFF; ram[1934] = 8'hFF; ram[1935] = 8'hFF;
        ram[1936] = 8'h0F; ram[1937] = 8'h0F; ram[1938] = 8'h0F; ram[1939] = 8'h00;
        ram[1940] = 8'h00; ram[1941] = 8'hFF; ram[1942] = 8'hFF; ram[1943] = 8'hFF;
        ram[1944] = 8'hFF; ram[1945] = 8'hFF; ram[1946] = 8'hFF; ram[1947] = 8'h00;
        ram[1948] = 8'h00; ram[1949] = 8'hFF; ram[1950] = 8'hFF; ram[1951] = 8'hFF;
        ram[1952] = 8'h00; ram[1953] = 8'h00; ram[1954] = 8'h00; ram[1955] = 8'hF0;
        ram[1956] = 8'hF0; ram[1957] = 8'hFF; ram[1958] = 8'hFF; ram[1959] = 8'hFF;
        ram[1960] = 8'hF0; ram[1961] = 8'hF0; ram[1962] = 8'hF0; ram[1963] = 8'hF0;
        ram[1964] = 8'hF0; ram[1965] = 8'hFF; ram[1966] = 8'hFF; ram[1967] = 8'hFF;
        ram[1968] = 8'h0F; ram[1969] = 8'h0F; ram[1970] = 8'h0F; ram[1971] = 8'hF0;
        ram[1972] = 8'hF0; ram[1973] = 8'hFF; ram[1974] = 8'hFF; ram[1975] = 8'hFF;
        ram[1976] = 8'hFF; ram[1977] = 8'hFF; ram[1978] = 8'hFF; ram[1979] = 8'hF0;
        ram[1980] = 8'hF0; ram[1981] = 8'hFF; ram[1982] = 8'hFF; ram[1983] = 8'hFF;
        ram[1984] = 8'h00; ram[1985] = 8'h00; ram[1986] = 8'h00; ram[1987] = 8'h0F;
        ram[1988] = 8'h0F; ram[1989] = 8'hFF; ram[1990] = 8'hFF; ram[1991] = 8'hFF;
        ram[1992] = 8'hF0; ram[1993] = 8'hF0; ram[1994] = 8'hF0; ram[1995] = 8'h0F;
        ram[1996] = 8'h0F; ram[1997] = 8'hFF; ram[1998] = 8'hFF; ram[1999] = 8'hFF;
        ram[2000] = 8'h0F; ram[2001] = 8'h0F; ram[2002] = 8'h0F; ram[2003] = 8'h0F;
        ram[2004] = 8'h0F; ram[2005] = 8'hFF; ram[2006] = 8'hFF; ram[2007] = 8'hFF;
        ram[2008] = 8'hFF; ram[2009] = 8'hFF; ram[2010] = 8'hFF; ram[2011] = 8'h0F;
        ram[2012] = 8'h0F; ram[2013] = 8'hFF; ram[2014] = 8'hFF; ram[2015] = 8'hFF;
        ram[2016] = 8'h00; ram[2017] = 8'h00; ram[2018] = 8'h00; ram[2019] = 8'hFF;
        ram[2020] = 8'hFF; ram[2021] = 8'hFF; ram[2022] = 8'hFF; ram[2023] = 8'hFF;
        ram[2024] = 8'hF0; ram[2025] = 8'hF0; ram[2026] = 8'hF0; ram[2027] = 8'hFF;
        ram[2028] = 8'hFF; ram[2029] = 8'hFF; ram[2030] = 8'hFF; ram[2031] = 8'hFF;
        ram[2032] = 8'h0F; ram[2033] = 8'h0F; ram[2034] = 8'h0F; ram[2035] = 8'hFF;
        ram[2036] = 8'hFF; ram[2037] = 8'hFF; ram[2038] = 8'hFF; ram[2039] = 8'hFF;
        ram[2040] = 8'hFF; ram[2041] = 8'hFF; ram[2042] = 8'hFF; ram[2043] = 8'hFF;
        ram[2044] = 8'hFF; ram[2045] = 8'hFF; ram[2046] = 8'hFF; ram[2047] = 8'hFF;
    end

    // always @(posedge clk)
    // begin
    //     if (wren1) ram[addr1] = wrdata1;
    //     rddata1 <= ram[addr1];
    // end

    always @(posedge clk)
    begin
        rddata2 <= ram[addr2];
    end

endmodule
