`timescale  1 ps / 1 ps


module BUFG (O, I);

    output O;

    input  I;


endmodule

