module bootrom(
    input  wire        clk,
    input  wire [12:0] addr,
    output reg   [7:0] rddata);

    always @(posedge(clk))
        case (addr)
            13'h0000: rddata <= 8'hC3;
            13'h0001: rddata <= 8'hE1;
            13'h0002: rddata <= 8'h1F;
            13'h0003: rddata <= 8'h82;
            13'h0004: rddata <= 8'h06;
            13'h0005: rddata <= 8'h22;
            13'h0006: rddata <= 8'h0B;
            13'h0007: rddata <= 8'h00;
            13'h0008: rddata <= 8'h7E;
            13'h0009: rddata <= 8'hE3;
            13'h000A: rddata <= 8'hBE;
            13'h000B: rddata <= 8'h23;
            13'h000C: rddata <= 8'hE3;
            13'h000D: rddata <= 8'hC2;
            13'h000E: rddata <= 8'hC4;
            13'h000F: rddata <= 8'h03;
            13'h0010: rddata <= 8'h23;
            13'h0011: rddata <= 8'h7E;
            13'h0012: rddata <= 8'hFE;
            13'h0013: rddata <= 8'h3A;
            13'h0014: rddata <= 8'hD0;
            13'h0015: rddata <= 8'hC3;
            13'h0016: rddata <= 8'h70;
            13'h0017: rddata <= 8'h06;
            13'h0018: rddata <= 8'hC3;
            13'h0019: rddata <= 8'h8A;
            13'h001A: rddata <= 8'h19;
            13'h001B: rddata <= 8'h00;
            13'h001C: rddata <= 8'h00;
            13'h001D: rddata <= 8'h00;
            13'h001E: rddata <= 8'h00;
            13'h001F: rddata <= 8'h00;
            13'h0020: rddata <= 8'h7C;
            13'h0021: rddata <= 8'h92;
            13'h0022: rddata <= 8'hC0;
            13'h0023: rddata <= 8'h7D;
            13'h0024: rddata <= 8'h93;
            13'h0025: rddata <= 8'hC9;
            13'h0026: rddata <= 8'h00;
            13'h0027: rddata <= 8'h00;
            13'h0028: rddata <= 8'h3A;
            13'h0029: rddata <= 8'hE7;
            13'h002A: rddata <= 8'h38;
            13'h002B: rddata <= 8'hB7;
            13'h002C: rddata <= 8'hC2;
            13'h002D: rddata <= 8'hEB;
            13'h002E: rddata <= 8'h14;
            13'h002F: rddata <= 8'hC9;
            13'h0030: rddata <= 8'hDD;
            13'h0031: rddata <= 8'h2A;
            13'h0032: rddata <= 8'h06;
            13'h0033: rddata <= 8'h38;
            13'h0034: rddata <= 8'hDD;
            13'h0035: rddata <= 8'hE9;
            13'h0036: rddata <= 8'h00;
            13'h0037: rddata <= 8'h00;
            13'h0038: rddata <= 8'hC3;
            13'h0039: rddata <= 8'h03;
            13'h003A: rddata <= 8'h38;
            13'h003B: rddata <= 8'hD9;
            13'h003C: rddata <= 8'hE1;
            13'h003D: rddata <= 8'h23;
            13'h003E: rddata <= 8'hE5;
            13'h003F: rddata <= 8'hD9;
            13'h0040: rddata <= 8'hC9;
            13'h0041: rddata <= 8'h31;
            13'h0042: rddata <= 8'hA0;
            13'h0043: rddata <= 8'h38;
            13'h0044: rddata <= 8'h3E;
            13'h0045: rddata <= 8'h0B;
            13'h0046: rddata <= 8'hCD;
            13'h0047: rddata <= 8'h94;
            13'h0048: rddata <= 8'h1D;
            13'h0049: rddata <= 8'h2A;
            13'h004A: rddata <= 8'h01;
            13'h004B: rddata <= 8'h38;
            13'h004C: rddata <= 8'h36;
            13'h004D: rddata <= 8'h20;
            13'h004E: rddata <= 8'h3E;
            13'h004F: rddata <= 8'h07;
            13'h0050: rddata <= 8'hCD;
            13'h0051: rddata <= 8'h94;
            13'h0052: rddata <= 8'h1D;
            13'h0053: rddata <= 8'hAF;
            13'h0054: rddata <= 8'hD3;
            13'h0055: rddata <= 8'hFF;
            13'h0056: rddata <= 8'h21;
            13'h0057: rddata <= 8'hFF;
            13'h0058: rddata <= 8'h2F;
            13'h0059: rddata <= 8'h22;
            13'h005A: rddata <= 8'h5D;
            13'h005B: rddata <= 8'h38;
            13'h005C: rddata <= 8'h11;
            13'h005D: rddata <= 8'h11;
            13'h005E: rddata <= 8'hE0;
            13'h005F: rddata <= 8'h21;
            13'h0060: rddata <= 8'h81;
            13'h0061: rddata <= 8'h00;
            13'h0062: rddata <= 8'h1B;
            13'h0063: rddata <= 8'h1B;
            13'h0064: rddata <= 8'h23;
            13'h0065: rddata <= 8'h1A;
            13'h0066: rddata <= 8'h0F;
            13'h0067: rddata <= 8'h0F;
            13'h0068: rddata <= 8'h83;
            13'h0069: rddata <= 8'hBE;
            13'h006A: rddata <= 8'h28;
            13'h006B: rddata <= 8'hF6;
            13'h006C: rddata <= 8'h7E;
            13'h006D: rddata <= 8'hB7;
            13'h006E: rddata <= 8'h20;
            13'h006F: rddata <= 8'h19;
            13'h0070: rddata <= 8'hEB;
            13'h0071: rddata <= 8'h06;
            13'h0072: rddata <= 8'h0C;
            13'h0073: rddata <= 8'h86;
            13'h0074: rddata <= 8'h23;
            13'h0075: rddata <= 8'h80;
            13'h0076: rddata <= 8'h05;
            13'h0077: rddata <= 8'h20;
            13'h0078: rddata <= 8'hFA;
            13'h0079: rddata <= 8'hAE;
            13'h007A: rddata <= 8'hD3;
            13'h007B: rddata <= 8'hFF;
            13'h007C: rddata <= 8'h32;
            13'h007D: rddata <= 8'h09;
            13'h007E: rddata <= 8'h38;
            13'h007F: rddata <= 8'hC3;
            13'h0080: rddata <= 8'h10;
            13'h0081: rddata <= 8'hE0;
            13'h0082: rddata <= 8'h2B;
            13'h0083: rddata <= 8'h37;
            13'h0084: rddata <= 8'h24;
            13'h0085: rddata <= 8'h24;
            13'h0086: rddata <= 8'h33;
            13'h0087: rddata <= 8'h2C;
            13'h0088: rddata <= 8'h00;
            13'h0089: rddata <= 8'h11;
            13'h008A: rddata <= 8'hA1;
            13'h008B: rddata <= 8'h31;
            13'h008C: rddata <= 8'h21;
            13'h008D: rddata <= 8'hB0;
            13'h008E: rddata <= 8'h00;
            13'h008F: rddata <= 8'h01;
            13'h0090: rddata <= 8'h05;
            13'h0091: rddata <= 8'h00;
            13'h0092: rddata <= 8'hED;
            13'h0093: rddata <= 8'hB0;
            13'h0094: rddata <= 8'h11;
            13'h0095: rddata <= 8'h10;
            13'h0096: rddata <= 8'h32;
            13'h0097: rddata <= 8'h21;
            13'h0098: rddata <= 8'hB5;
            13'h0099: rddata <= 8'h00;
            13'h009A: rddata <= 8'h01;
            13'h009B: rddata <= 8'h19;
            13'h009C: rddata <= 8'h00;
            13'h009D: rddata <= 8'hED;
            13'h009E: rddata <= 8'hB0;
            13'h009F: rddata <= 8'h06;
            13'h00A0: rddata <= 8'h03;
            13'h00A1: rddata <= 8'hCD;
            13'h00A2: rddata <= 8'hCF;
            13'h00A3: rddata <= 8'h00;
            13'h00A4: rddata <= 8'h06;
            13'h00A5: rddata <= 8'h02;
            13'h00A6: rddata <= 8'hCD;
            13'h00A7: rddata <= 8'hCF;
            13'h00A8: rddata <= 8'h00;
            13'h00A9: rddata <= 8'h06;
            13'h00AA: rddata <= 8'h06;
            13'h00AB: rddata <= 8'hCD;
            13'h00AC: rddata <= 8'hCF;
            13'h00AD: rddata <= 8'h00;
            13'h00AE: rddata <= 8'h18;
            13'h00AF: rddata <= 8'hEF;
            13'h00B0: rddata <= 8'h42;
            13'h00B1: rddata <= 8'h41;
            13'h00B2: rddata <= 8'h53;
            13'h00B3: rddata <= 8'h49;
            13'h00B4: rddata <= 8'h43;
            13'h00B5: rddata <= 8'h50;
            13'h00B6: rddata <= 8'h72;
            13'h00B7: rddata <= 8'h65;
            13'h00B8: rddata <= 8'h73;
            13'h00B9: rddata <= 8'h73;
            13'h00BA: rddata <= 8'h20;
            13'h00BB: rddata <= 8'h52;
            13'h00BC: rddata <= 8'h45;
            13'h00BD: rddata <= 8'h54;
            13'h00BE: rddata <= 8'h55;
            13'h00BF: rddata <= 8'h52;
            13'h00C0: rddata <= 8'h4E;
            13'h00C1: rddata <= 8'h20;
            13'h00C2: rddata <= 8'h6B;
            13'h00C3: rddata <= 8'h65;
            13'h00C4: rddata <= 8'h79;
            13'h00C5: rddata <= 8'h20;
            13'h00C6: rddata <= 8'h74;
            13'h00C7: rddata <= 8'h6F;
            13'h00C8: rddata <= 8'h20;
            13'h00C9: rddata <= 8'h73;
            13'h00CA: rddata <= 8'h74;
            13'h00CB: rddata <= 8'h61;
            13'h00CC: rddata <= 8'h72;
            13'h00CD: rddata <= 8'h74;
            13'h00CE: rddata <= 8'h00;
            13'h00CF: rddata <= 8'h21;
            13'h00D0: rddata <= 8'h00;
            13'h00D1: rddata <= 8'h34;
            13'h00D2: rddata <= 8'h70;
            13'h00D3: rddata <= 8'h23;
            13'h00D4: rddata <= 8'h7C;
            13'h00D5: rddata <= 8'hFE;
            13'h00D6: rddata <= 8'h38;
            13'h00D7: rddata <= 8'h20;
            13'h00D8: rddata <= 8'hF9;
            13'h00D9: rddata <= 8'h21;
            13'h00DA: rddata <= 8'h00;
            13'h00DB: rddata <= 8'h40;
            13'h00DC: rddata <= 8'hCD;
            13'h00DD: rddata <= 8'h80;
            13'h00DE: rddata <= 8'h1E;
            13'h00DF: rddata <= 8'hFE;
            13'h00E0: rddata <= 8'h0D;
            13'h00E1: rddata <= 8'h28;
            13'h00E2: rddata <= 8'h1A;
            13'h00E3: rddata <= 8'hFE;
            13'h00E4: rddata <= 8'h03;
            13'h00E5: rddata <= 8'h28;
            13'h00E6: rddata <= 8'h06;
            13'h00E7: rddata <= 8'h2B;
            13'h00E8: rddata <= 8'h7C;
            13'h00E9: rddata <= 8'hB5;
            13'h00EA: rddata <= 8'h20;
            13'h00EB: rddata <= 8'hF0;
            13'h00EC: rddata <= 8'hC9;
            13'h00ED: rddata <= 8'h3E;
            13'h00EE: rddata <= 8'h0B;
            13'h00EF: rddata <= 8'hCD;
            13'h00F0: rddata <= 8'h72;
            13'h00F1: rddata <= 8'h1D;
            13'h00F2: rddata <= 8'h3A;
            13'h00F3: rddata <= 8'h09;
            13'h00F4: rddata <= 8'h38;
            13'h00F5: rddata <= 8'hD3;
            13'h00F6: rddata <= 8'hFF;
            13'h00F7: rddata <= 8'hCD;
            13'h00F8: rddata <= 8'hE5;
            13'h00F9: rddata <= 8'h0B;
            13'h00FA: rddata <= 8'hCD;
            13'h00FB: rddata <= 8'h40;
            13'h00FC: rddata <= 8'h1A;
            13'h00FD: rddata <= 8'h21;
            13'h00FE: rddata <= 8'h87;
            13'h00FF: rddata <= 8'h01;
            13'h0100: rddata <= 8'h01;
            13'h0101: rddata <= 8'h51;
            13'h0102: rddata <= 8'h00;
            13'h0103: rddata <= 8'h11;
            13'h0104: rddata <= 8'h03;
            13'h0105: rddata <= 8'h38;
            13'h0106: rddata <= 8'hED;
            13'h0107: rddata <= 8'hB0;
            13'h0108: rddata <= 8'hAF;
            13'h0109: rddata <= 8'h32;
            13'h010A: rddata <= 8'hA9;
            13'h010B: rddata <= 8'h38;
            13'h010C: rddata <= 8'h32;
            13'h010D: rddata <= 8'h00;
            13'h010E: rddata <= 8'h39;
            13'h010F: rddata <= 8'h21;
            13'h0110: rddata <= 8'h64;
            13'h0111: rddata <= 8'h39;
            13'h0112: rddata <= 8'h23;
            13'h0113: rddata <= 8'h4E;
            13'h0114: rddata <= 8'h7C;
            13'h0115: rddata <= 8'hB5;
            13'h0116: rddata <= 8'h28;
            13'h0117: rddata <= 8'h0B;
            13'h0118: rddata <= 8'hA9;
            13'h0119: rddata <= 8'h77;
            13'h011A: rddata <= 8'h46;
            13'h011B: rddata <= 8'h2F;
            13'h011C: rddata <= 8'h77;
            13'h011D: rddata <= 8'h7E;
            13'h011E: rddata <= 8'h2F;
            13'h011F: rddata <= 8'h71;
            13'h0120: rddata <= 8'hB8;
            13'h0121: rddata <= 8'h28;
            13'h0122: rddata <= 8'hEF;
            13'h0123: rddata <= 8'h2B;
            13'h0124: rddata <= 8'h11;
            13'h0125: rddata <= 8'h2C;
            13'h0126: rddata <= 8'h3A;
            13'h0127: rddata <= 8'hE7;
            13'h0128: rddata <= 8'hDA;
            13'h0129: rddata <= 8'hB7;
            13'h012A: rddata <= 8'h0B;
            13'h012B: rddata <= 8'h11;
            13'h012C: rddata <= 8'hCE;
            13'h012D: rddata <= 8'hFF;
            13'h012E: rddata <= 8'h22;
            13'h012F: rddata <= 8'hAD;
            13'h0130: rddata <= 8'h38;
            13'h0131: rddata <= 8'h19;
            13'h0132: rddata <= 8'h22;
            13'h0133: rddata <= 8'h4B;
            13'h0134: rddata <= 8'h38;
            13'h0135: rddata <= 8'hCD;
            13'h0136: rddata <= 8'hBE;
            13'h0137: rddata <= 8'h0B;
            13'h0138: rddata <= 8'hCD;
            13'h0139: rddata <= 8'hF2;
            13'h013A: rddata <= 8'h1F;
            13'h013B: rddata <= 8'h31;
            13'h013C: rddata <= 8'h65;
            13'h013D: rddata <= 8'h38;
            13'h013E: rddata <= 8'hCD;
            13'h013F: rddata <= 8'hE5;
            13'h0140: rddata <= 8'h0B;
            13'h0141: rddata <= 8'h21;
            13'h0142: rddata <= 8'h05;
            13'h0143: rddata <= 8'h20;
            13'h0144: rddata <= 8'h11;
            13'h0145: rddata <= 8'h82;
            13'h0146: rddata <= 8'h00;
            13'h0147: rddata <= 8'h1A;
            13'h0148: rddata <= 8'hB7;
            13'h0149: rddata <= 8'hCA;
            13'h014A: rddata <= 8'hE8;
            13'h014B: rddata <= 8'h1F;
            13'h014C: rddata <= 8'hBE;
            13'h014D: rddata <= 8'h20;
            13'h014E: rddata <= 8'h04;
            13'h014F: rddata <= 8'h2B;
            13'h0150: rddata <= 8'h13;
            13'h0151: rddata <= 8'h18;
            13'h0152: rddata <= 8'hF4;
            13'h0153: rddata <= 8'hED;
            13'h0154: rddata <= 8'h5F;
            13'h0155: rddata <= 8'h17;
            13'h0156: rddata <= 8'h81;
            13'h0157: rddata <= 8'hD3;
            13'h0158: rddata <= 8'hFF;
            13'h0159: rddata <= 8'h32;
            13'h015A: rddata <= 8'h09;
            13'h015B: rddata <= 8'h38;
            13'h015C: rddata <= 8'hC3;
            13'h015D: rddata <= 8'h02;
            13'h015E: rddata <= 8'h04;
            13'h015F: rddata <= 8'h0B;
            13'h0160: rddata <= 8'h43;
            13'h0161: rddata <= 8'h6F;
            13'h0162: rddata <= 8'h70;
            13'h0163: rddata <= 8'h79;
            13'h0164: rddata <= 8'h72;
            13'h0165: rddata <= 8'h69;
            13'h0166: rddata <= 8'h67;
            13'h0167: rddata <= 8'h68;
            13'h0168: rddata <= 8'h74;
            13'h0169: rddata <= 8'h20;
            13'h016A: rddata <= 8'h05;
            13'h016B: rddata <= 8'h20;
            13'h016C: rddata <= 8'h31;
            13'h016D: rddata <= 8'h39;
            13'h016E: rddata <= 8'h38;
            13'h016F: rddata <= 8'h32;
            13'h0170: rddata <= 8'h20;
            13'h0171: rddata <= 8'h62;
            13'h0172: rddata <= 8'h79;
            13'h0173: rddata <= 8'h20;
            13'h0174: rddata <= 8'h4D;
            13'h0175: rddata <= 8'h69;
            13'h0176: rddata <= 8'h63;
            13'h0177: rddata <= 8'h72;
            13'h0178: rddata <= 8'h6F;
            13'h0179: rddata <= 8'h73;
            13'h017A: rddata <= 8'h6F;
            13'h017B: rddata <= 8'h66;
            13'h017C: rddata <= 8'h74;
            13'h017D: rddata <= 8'h20;
            13'h017E: rddata <= 8'h49;
            13'h017F: rddata <= 8'h6E;
            13'h0180: rddata <= 8'h63;
            13'h0181: rddata <= 8'h2E;
            13'h0182: rddata <= 8'h20;
            13'h0183: rddata <= 8'h53;
            13'h0184: rddata <= 8'h32;
            13'h0185: rddata <= 8'h0A;
            13'h0186: rddata <= 8'h00;
            13'h0187: rddata <= 8'hC3;
            13'h0188: rddata <= 8'h97;
            13'h0189: rddata <= 8'h06;
            13'h018A: rddata <= 8'h3B;
            13'h018B: rddata <= 8'h00;
            13'h018C: rddata <= 8'h00;
            13'h018D: rddata <= 8'hA3;
            13'h018E: rddata <= 8'h00;
            13'h018F: rddata <= 8'h00;
            13'h0190: rddata <= 8'h00;
            13'h0191: rddata <= 8'h20;
            13'h0192: rddata <= 8'h00;
            13'h0193: rddata <= 8'h00;
            13'h0194: rddata <= 8'hD6;
            13'h0195: rddata <= 8'h00;
            13'h0196: rddata <= 8'h6F;
            13'h0197: rddata <= 8'h7C;
            13'h0198: rddata <= 8'hDE;
            13'h0199: rddata <= 8'h00;
            13'h019A: rddata <= 8'h67;
            13'h019B: rddata <= 8'h78;
            13'h019C: rddata <= 8'hDE;
            13'h019D: rddata <= 8'h00;
            13'h019E: rddata <= 8'h47;
            13'h019F: rddata <= 8'h3E;
            13'h01A0: rddata <= 8'h00;
            13'h01A1: rddata <= 8'hC9;
            13'h01A2: rddata <= 8'h00;
            13'h01A3: rddata <= 8'h00;
            13'h01A4: rddata <= 8'h00;
            13'h01A5: rddata <= 8'h35;
            13'h01A6: rddata <= 8'h4A;
            13'h01A7: rddata <= 8'hCA;
            13'h01A8: rddata <= 8'h99;
            13'h01A9: rddata <= 8'h39;
            13'h01AA: rddata <= 8'h1C;
            13'h01AB: rddata <= 8'h76;
            13'h01AC: rddata <= 8'h98;
            13'h01AD: rddata <= 8'h22;
            13'h01AE: rddata <= 8'h95;
            13'h01AF: rddata <= 8'hB3;
            13'h01B0: rddata <= 8'h98;
            13'h01B1: rddata <= 8'h0A;
            13'h01B2: rddata <= 8'hDD;
            13'h01B3: rddata <= 8'h47;
            13'h01B4: rddata <= 8'h98;
            13'h01B5: rddata <= 8'h53;
            13'h01B6: rddata <= 8'hD1;
            13'h01B7: rddata <= 8'h99;
            13'h01B8: rddata <= 8'h99;
            13'h01B9: rddata <= 8'h0A;
            13'h01BA: rddata <= 8'h1A;
            13'h01BB: rddata <= 8'h9F;
            13'h01BC: rddata <= 8'h98;
            13'h01BD: rddata <= 8'h65;
            13'h01BE: rddata <= 8'hBC;
            13'h01BF: rddata <= 8'hCD;
            13'h01C0: rddata <= 8'h98;
            13'h01C1: rddata <= 8'hD6;
            13'h01C2: rddata <= 8'h77;
            13'h01C3: rddata <= 8'h3E;
            13'h01C4: rddata <= 8'h98;
            13'h01C5: rddata <= 8'h52;
            13'h01C6: rddata <= 8'hC7;
            13'h01C7: rddata <= 8'h4F;
            13'h01C8: rddata <= 8'h80;
            13'h01C9: rddata <= 8'h00;
            13'h01CA: rddata <= 8'h00;
            13'h01CB: rddata <= 8'h00;
            13'h01CC: rddata <= 8'h28;
            13'h01CD: rddata <= 8'h0E;
            13'h01CE: rddata <= 8'h00;
            13'h01CF: rddata <= 8'h64;
            13'h01D0: rddata <= 8'h39;
            13'h01D1: rddata <= 8'hFE;
            13'h01D2: rddata <= 8'hFF;
            13'h01D3: rddata <= 8'h01;
            13'h01D4: rddata <= 8'h39;
            13'h01D5: rddata <= 8'h21;
            13'h01D6: rddata <= 8'h0C;
            13'h01D7: rddata <= 8'hBC;
            13'h01D8: rddata <= 8'h05;
            13'h01D9: rddata <= 8'h13;
            13'h01DA: rddata <= 8'h0D;
            13'h01DB: rddata <= 8'h1C;
            13'h01DC: rddata <= 8'h07;
            13'h01DD: rddata <= 8'h93;
            13'h01DE: rddata <= 8'h08;
            13'h01DF: rddata <= 8'hCC;
            13'h01E0: rddata <= 8'h10;
            13'h01E1: rddata <= 8'hBE;
            13'h01E2: rddata <= 8'h08;
            13'h01E3: rddata <= 8'h31;
            13'h01E4: rddata <= 8'h07;
            13'h01E5: rddata <= 8'hDC;
            13'h01E6: rddata <= 8'h06;
            13'h01E7: rddata <= 8'hBE;
            13'h01E8: rddata <= 8'h06;
            13'h01E9: rddata <= 8'h9C;
            13'h01EA: rddata <= 8'h07;
            13'h01EB: rddata <= 8'h05;
            13'h01EC: rddata <= 8'h0C;
            13'h01ED: rddata <= 8'hCB;
            13'h01EE: rddata <= 8'h06;
            13'h01EF: rddata <= 8'hF8;
            13'h01F0: rddata <= 8'h06;
            13'h01F1: rddata <= 8'h1E;
            13'h01F2: rddata <= 8'h07;
            13'h01F3: rddata <= 8'h1F;
            13'h01F4: rddata <= 8'h0C;
            13'h01F5: rddata <= 8'h80;
            13'h01F6: rddata <= 8'h07;
            13'h01F7: rddata <= 8'hB5;
            13'h01F8: rddata <= 8'h07;
            13'h01F9: rddata <= 8'h15;
            13'h01FA: rddata <= 8'h1B;
            13'h01FB: rddata <= 8'h3B;
            13'h01FC: rddata <= 8'h0B;
            13'h01FD: rddata <= 8'h6D;
            13'h01FE: rddata <= 8'h0B;
            13'h01FF: rddata <= 8'hBC;
            13'h0200: rddata <= 8'h07;
            13'h0201: rddata <= 8'h4B;
            13'h0202: rddata <= 8'h0C;
            13'h0203: rddata <= 8'h6C;
            13'h0204: rddata <= 8'h05;
            13'h0205: rddata <= 8'h67;
            13'h0206: rddata <= 8'h05;
            13'h0207: rddata <= 8'hCD;
            13'h0208: rddata <= 8'h0C;
            13'h0209: rddata <= 8'h2C;
            13'h020A: rddata <= 8'h1C;
            13'h020B: rddata <= 8'h08;
            13'h020C: rddata <= 8'h1C;
            13'h020D: rddata <= 8'h4F;
            13'h020E: rddata <= 8'h1A;
            13'h020F: rddata <= 8'h4C;
            13'h0210: rddata <= 8'h1A;
            13'h0211: rddata <= 8'hD6;
            13'h0212: rddata <= 8'h1A;
            13'h0213: rddata <= 8'hBD;
            13'h0214: rddata <= 8'h0B;
            13'h0215: rddata <= 8'hF5;
            13'h0216: rddata <= 8'h14;
            13'h0217: rddata <= 8'hB1;
            13'h0218: rddata <= 8'h15;
            13'h0219: rddata <= 8'h09;
            13'h021A: rddata <= 8'h15;
            13'h021B: rddata <= 8'h03;
            13'h021C: rddata <= 8'h38;
            13'h021D: rddata <= 8'hA8;
            13'h021E: rddata <= 8'h10;
            13'h021F: rddata <= 8'h2E;
            13'h0220: rddata <= 8'h0B;
            13'h0221: rddata <= 8'h33;
            13'h0222: rddata <= 8'h0B;
            13'h0223: rddata <= 8'h75;
            13'h0224: rddata <= 8'h17;
            13'h0225: rddata <= 8'h66;
            13'h0226: rddata <= 8'h18;
            13'h0227: rddata <= 8'h85;
            13'h0228: rddata <= 8'h13;
            13'h0229: rddata <= 8'hCD;
            13'h022A: rddata <= 8'h17;
            13'h022B: rddata <= 8'hD7;
            13'h022C: rddata <= 8'h18;
            13'h022D: rddata <= 8'hDD;
            13'h022E: rddata <= 8'h18;
            13'h022F: rddata <= 8'h70;
            13'h0230: rddata <= 8'h19;
            13'h0231: rddata <= 8'h85;
            13'h0232: rddata <= 8'h19;
            13'h0233: rddata <= 8'h63;
            13'h0234: rddata <= 8'h0B;
            13'h0235: rddata <= 8'hF3;
            13'h0236: rddata <= 8'h0F;
            13'h0237: rddata <= 8'h29;
            13'h0238: rddata <= 8'h0E;
            13'h0239: rddata <= 8'h84;
            13'h023A: rddata <= 8'h10;
            13'h023B: rddata <= 8'h02;
            13'h023C: rddata <= 8'h10;
            13'h023D: rddata <= 8'h13;
            13'h023E: rddata <= 8'h10;
            13'h023F: rddata <= 8'h21;
            13'h0240: rddata <= 8'h10;
            13'h0241: rddata <= 8'h50;
            13'h0242: rddata <= 8'h10;
            13'h0243: rddata <= 8'h59;
            13'h0244: rddata <= 8'h10;
            13'h0245: rddata <= 8'hC5;
            13'h0246: rddata <= 8'h4E;
            13'h0247: rddata <= 8'h44;
            13'h0248: rddata <= 8'hC6;
            13'h0249: rddata <= 8'h4F;
            13'h024A: rddata <= 8'h52;
            13'h024B: rddata <= 8'hCE;
            13'h024C: rddata <= 8'h45;
            13'h024D: rddata <= 8'h58;
            13'h024E: rddata <= 8'h54;
            13'h024F: rddata <= 8'hC4;
            13'h0250: rddata <= 8'h41;
            13'h0251: rddata <= 8'h54;
            13'h0252: rddata <= 8'h41;
            13'h0253: rddata <= 8'hC9;
            13'h0254: rddata <= 8'h4E;
            13'h0255: rddata <= 8'h50;
            13'h0256: rddata <= 8'h55;
            13'h0257: rddata <= 8'h54;
            13'h0258: rddata <= 8'hC4;
            13'h0259: rddata <= 8'h49;
            13'h025A: rddata <= 8'h4D;
            13'h025B: rddata <= 8'hD2;
            13'h025C: rddata <= 8'h45;
            13'h025D: rddata <= 8'h41;
            13'h025E: rddata <= 8'h44;
            13'h025F: rddata <= 8'hCC;
            13'h0260: rddata <= 8'h45;
            13'h0261: rddata <= 8'h54;
            13'h0262: rddata <= 8'hC7;
            13'h0263: rddata <= 8'h4F;
            13'h0264: rddata <= 8'h54;
            13'h0265: rddata <= 8'h4F;
            13'h0266: rddata <= 8'hD2;
            13'h0267: rddata <= 8'h55;
            13'h0268: rddata <= 8'h4E;
            13'h0269: rddata <= 8'hC9;
            13'h026A: rddata <= 8'h46;
            13'h026B: rddata <= 8'hD2;
            13'h026C: rddata <= 8'h45;
            13'h026D: rddata <= 8'h53;
            13'h026E: rddata <= 8'h54;
            13'h026F: rddata <= 8'h4F;
            13'h0270: rddata <= 8'h52;
            13'h0271: rddata <= 8'h45;
            13'h0272: rddata <= 8'hC7;
            13'h0273: rddata <= 8'h4F;
            13'h0274: rddata <= 8'h53;
            13'h0275: rddata <= 8'h55;
            13'h0276: rddata <= 8'h42;
            13'h0277: rddata <= 8'hD2;
            13'h0278: rddata <= 8'h45;
            13'h0279: rddata <= 8'h54;
            13'h027A: rddata <= 8'h55;
            13'h027B: rddata <= 8'h52;
            13'h027C: rddata <= 8'h4E;
            13'h027D: rddata <= 8'hD2;
            13'h027E: rddata <= 8'h45;
            13'h027F: rddata <= 8'h4D;
            13'h0280: rddata <= 8'hD3;
            13'h0281: rddata <= 8'h54;
            13'h0282: rddata <= 8'h4F;
            13'h0283: rddata <= 8'h50;
            13'h0284: rddata <= 8'hCF;
            13'h0285: rddata <= 8'h4E;
            13'h0286: rddata <= 8'hCC;
            13'h0287: rddata <= 8'h50;
            13'h0288: rddata <= 8'h52;
            13'h0289: rddata <= 8'h49;
            13'h028A: rddata <= 8'h4E;
            13'h028B: rddata <= 8'h54;
            13'h028C: rddata <= 8'hC3;
            13'h028D: rddata <= 8'h4F;
            13'h028E: rddata <= 8'h50;
            13'h028F: rddata <= 8'h59;
            13'h0290: rddata <= 8'hC4;
            13'h0291: rddata <= 8'h45;
            13'h0292: rddata <= 8'h46;
            13'h0293: rddata <= 8'hD0;
            13'h0294: rddata <= 8'h4F;
            13'h0295: rddata <= 8'h4B;
            13'h0296: rddata <= 8'h45;
            13'h0297: rddata <= 8'hD0;
            13'h0298: rddata <= 8'h52;
            13'h0299: rddata <= 8'h49;
            13'h029A: rddata <= 8'h4E;
            13'h029B: rddata <= 8'h54;
            13'h029C: rddata <= 8'hC3;
            13'h029D: rddata <= 8'h4F;
            13'h029E: rddata <= 8'h4E;
            13'h029F: rddata <= 8'h54;
            13'h02A0: rddata <= 8'hCC;
            13'h02A1: rddata <= 8'h49;
            13'h02A2: rddata <= 8'h53;
            13'h02A3: rddata <= 8'h54;
            13'h02A4: rddata <= 8'hCC;
            13'h02A5: rddata <= 8'h4C;
            13'h02A6: rddata <= 8'h49;
            13'h02A7: rddata <= 8'h53;
            13'h02A8: rddata <= 8'h54;
            13'h02A9: rddata <= 8'hC3;
            13'h02AA: rddata <= 8'h4C;
            13'h02AB: rddata <= 8'h45;
            13'h02AC: rddata <= 8'h41;
            13'h02AD: rddata <= 8'h52;
            13'h02AE: rddata <= 8'hC3;
            13'h02AF: rddata <= 8'h4C;
            13'h02B0: rddata <= 8'h4F;
            13'h02B1: rddata <= 8'h41;
            13'h02B2: rddata <= 8'h44;
            13'h02B3: rddata <= 8'hC3;
            13'h02B4: rddata <= 8'h53;
            13'h02B5: rddata <= 8'h41;
            13'h02B6: rddata <= 8'h56;
            13'h02B7: rddata <= 8'h45;
            13'h02B8: rddata <= 8'hD0;
            13'h02B9: rddata <= 8'h53;
            13'h02BA: rddata <= 8'h45;
            13'h02BB: rddata <= 8'h54;
            13'h02BC: rddata <= 8'hD0;
            13'h02BD: rddata <= 8'h52;
            13'h02BE: rddata <= 8'h45;
            13'h02BF: rddata <= 8'h53;
            13'h02C0: rddata <= 8'h45;
            13'h02C1: rddata <= 8'h54;
            13'h02C2: rddata <= 8'hD3;
            13'h02C3: rddata <= 8'h4F;
            13'h02C4: rddata <= 8'h55;
            13'h02C5: rddata <= 8'h4E;
            13'h02C6: rddata <= 8'h44;
            13'h02C7: rddata <= 8'hCE;
            13'h02C8: rddata <= 8'h45;
            13'h02C9: rddata <= 8'h57;
            13'h02CA: rddata <= 8'hD4;
            13'h02CB: rddata <= 8'h41;
            13'h02CC: rddata <= 8'h42;
            13'h02CD: rddata <= 8'h28;
            13'h02CE: rddata <= 8'hD4;
            13'h02CF: rddata <= 8'h4F;
            13'h02D0: rddata <= 8'hC6;
            13'h02D1: rddata <= 8'h4E;
            13'h02D2: rddata <= 8'hD3;
            13'h02D3: rddata <= 8'h50;
            13'h02D4: rddata <= 8'h43;
            13'h02D5: rddata <= 8'h28;
            13'h02D6: rddata <= 8'hC9;
            13'h02D7: rddata <= 8'h4E;
            13'h02D8: rddata <= 8'h4B;
            13'h02D9: rddata <= 8'h45;
            13'h02DA: rddata <= 8'h59;
            13'h02DB: rddata <= 8'h24;
            13'h02DC: rddata <= 8'hD4;
            13'h02DD: rddata <= 8'h48;
            13'h02DE: rddata <= 8'h45;
            13'h02DF: rddata <= 8'h4E;
            13'h02E0: rddata <= 8'hCE;
            13'h02E1: rddata <= 8'h4F;
            13'h02E2: rddata <= 8'h54;
            13'h02E3: rddata <= 8'hD3;
            13'h02E4: rddata <= 8'h54;
            13'h02E5: rddata <= 8'h45;
            13'h02E6: rddata <= 8'h50;
            13'h02E7: rddata <= 8'hAB;
            13'h02E8: rddata <= 8'hAD;
            13'h02E9: rddata <= 8'hAA;
            13'h02EA: rddata <= 8'hAF;
            13'h02EB: rddata <= 8'hDE;
            13'h02EC: rddata <= 8'hC1;
            13'h02ED: rddata <= 8'h4E;
            13'h02EE: rddata <= 8'h44;
            13'h02EF: rddata <= 8'hCF;
            13'h02F0: rddata <= 8'h52;
            13'h02F1: rddata <= 8'hBE;
            13'h02F2: rddata <= 8'hBD;
            13'h02F3: rddata <= 8'hBC;
            13'h02F4: rddata <= 8'hD3;
            13'h02F5: rddata <= 8'h47;
            13'h02F6: rddata <= 8'h4E;
            13'h02F7: rddata <= 8'hC9;
            13'h02F8: rddata <= 8'h4E;
            13'h02F9: rddata <= 8'h54;
            13'h02FA: rddata <= 8'hC1;
            13'h02FB: rddata <= 8'h42;
            13'h02FC: rddata <= 8'h53;
            13'h02FD: rddata <= 8'hD5;
            13'h02FE: rddata <= 8'h53;
            13'h02FF: rddata <= 8'h52;
            13'h0300: rddata <= 8'hC6;
            13'h0301: rddata <= 8'h52;
            13'h0302: rddata <= 8'h45;
            13'h0303: rddata <= 8'hCC;
            13'h0304: rddata <= 8'h50;
            13'h0305: rddata <= 8'h4F;
            13'h0306: rddata <= 8'h53;
            13'h0307: rddata <= 8'hD0;
            13'h0308: rddata <= 8'h4F;
            13'h0309: rddata <= 8'h53;
            13'h030A: rddata <= 8'hD3;
            13'h030B: rddata <= 8'h51;
            13'h030C: rddata <= 8'h52;
            13'h030D: rddata <= 8'hD2;
            13'h030E: rddata <= 8'h4E;
            13'h030F: rddata <= 8'h44;
            13'h0310: rddata <= 8'hCC;
            13'h0311: rddata <= 8'h4F;
            13'h0312: rddata <= 8'h47;
            13'h0313: rddata <= 8'hC5;
            13'h0314: rddata <= 8'h58;
            13'h0315: rddata <= 8'h50;
            13'h0316: rddata <= 8'hC3;
            13'h0317: rddata <= 8'h4F;
            13'h0318: rddata <= 8'h53;
            13'h0319: rddata <= 8'hD3;
            13'h031A: rddata <= 8'h49;
            13'h031B: rddata <= 8'h4E;
            13'h031C: rddata <= 8'hD4;
            13'h031D: rddata <= 8'h41;
            13'h031E: rddata <= 8'h4E;
            13'h031F: rddata <= 8'hC1;
            13'h0320: rddata <= 8'h54;
            13'h0321: rddata <= 8'h4E;
            13'h0322: rddata <= 8'hD0;
            13'h0323: rddata <= 8'h45;
            13'h0324: rddata <= 8'h45;
            13'h0325: rddata <= 8'h4B;
            13'h0326: rddata <= 8'hCC;
            13'h0327: rddata <= 8'h45;
            13'h0328: rddata <= 8'h4E;
            13'h0329: rddata <= 8'hD3;
            13'h032A: rddata <= 8'h54;
            13'h032B: rddata <= 8'h52;
            13'h032C: rddata <= 8'h24;
            13'h032D: rddata <= 8'hD6;
            13'h032E: rddata <= 8'h41;
            13'h032F: rddata <= 8'h4C;
            13'h0330: rddata <= 8'hC1;
            13'h0331: rddata <= 8'h53;
            13'h0332: rddata <= 8'h43;
            13'h0333: rddata <= 8'hC3;
            13'h0334: rddata <= 8'h48;
            13'h0335: rddata <= 8'h52;
            13'h0336: rddata <= 8'h24;
            13'h0337: rddata <= 8'hCC;
            13'h0338: rddata <= 8'h45;
            13'h0339: rddata <= 8'h46;
            13'h033A: rddata <= 8'h54;
            13'h033B: rddata <= 8'h24;
            13'h033C: rddata <= 8'hD2;
            13'h033D: rddata <= 8'h49;
            13'h033E: rddata <= 8'h47;
            13'h033F: rddata <= 8'h48;
            13'h0340: rddata <= 8'h54;
            13'h0341: rddata <= 8'h24;
            13'h0342: rddata <= 8'hCD;
            13'h0343: rddata <= 8'h49;
            13'h0344: rddata <= 8'h44;
            13'h0345: rddata <= 8'h24;
            13'h0346: rddata <= 8'hD0;
            13'h0347: rddata <= 8'h4F;
            13'h0348: rddata <= 8'h49;
            13'h0349: rddata <= 8'h4E;
            13'h034A: rddata <= 8'h54;
            13'h034B: rddata <= 8'h80;
            13'h034C: rddata <= 8'h79;
            13'h034D: rddata <= 8'h5C;
            13'h034E: rddata <= 8'h16;
            13'h034F: rddata <= 8'h79;
            13'h0350: rddata <= 8'h5C;
            13'h0351: rddata <= 8'h12;
            13'h0352: rddata <= 8'h7C;
            13'h0353: rddata <= 8'hC9;
            13'h0354: rddata <= 8'h13;
            13'h0355: rddata <= 8'h7C;
            13'h0356: rddata <= 8'h2D;
            13'h0357: rddata <= 8'h14;
            13'h0358: rddata <= 8'h7F;
            13'h0359: rddata <= 8'h7E;
            13'h035A: rddata <= 8'h17;
            13'h035B: rddata <= 8'h50;
            13'h035C: rddata <= 8'hA9;
            13'h035D: rddata <= 8'h0A;
            13'h035E: rddata <= 8'h46;
            13'h035F: rddata <= 8'hA8;
            13'h0360: rddata <= 8'h0A;
            13'h0361: rddata <= 8'h20;
            13'h0362: rddata <= 8'h45;
            13'h0363: rddata <= 8'h72;
            13'h0364: rddata <= 8'h72;
            13'h0365: rddata <= 8'h6F;
            13'h0366: rddata <= 8'h72;
            13'h0367: rddata <= 8'h07;
            13'h0368: rddata <= 8'h00;
            13'h0369: rddata <= 8'h20;
            13'h036A: rddata <= 8'h69;
            13'h036B: rddata <= 8'h6E;
            13'h036C: rddata <= 8'h20;
            13'h036D: rddata <= 8'h00;
            13'h036E: rddata <= 8'h4F;
            13'h036F: rddata <= 8'h6B;
            13'h0370: rddata <= 8'h0D;
            13'h0371: rddata <= 8'h0A;
            13'h0372: rddata <= 8'h00;
            13'h0373: rddata <= 8'h42;
            13'h0374: rddata <= 8'h72;
            13'h0375: rddata <= 8'h65;
            13'h0376: rddata <= 8'h61;
            13'h0377: rddata <= 8'h6B;
            13'h0378: rddata <= 8'h00;
            13'h0379: rddata <= 8'h4E;
            13'h037A: rddata <= 8'h46;
            13'h037B: rddata <= 8'h53;
            13'h037C: rddata <= 8'h4E;
            13'h037D: rddata <= 8'h52;
            13'h037E: rddata <= 8'h47;
            13'h037F: rddata <= 8'h4F;
            13'h0380: rddata <= 8'h44;
            13'h0381: rddata <= 8'h46;
            13'h0382: rddata <= 8'h43;
            13'h0383: rddata <= 8'h4F;
            13'h0384: rddata <= 8'h56;
            13'h0385: rddata <= 8'h4F;
            13'h0386: rddata <= 8'h4D;
            13'h0387: rddata <= 8'h55;
            13'h0388: rddata <= 8'h4C;
            13'h0389: rddata <= 8'h42;
            13'h038A: rddata <= 8'h53;
            13'h038B: rddata <= 8'h44;
            13'h038C: rddata <= 8'h44;
            13'h038D: rddata <= 8'h2F;
            13'h038E: rddata <= 8'h30;
            13'h038F: rddata <= 8'h49;
            13'h0390: rddata <= 8'h44;
            13'h0391: rddata <= 8'h54;
            13'h0392: rddata <= 8'h4D;
            13'h0393: rddata <= 8'h4F;
            13'h0394: rddata <= 8'h53;
            13'h0395: rddata <= 8'h4C;
            13'h0396: rddata <= 8'h53;
            13'h0397: rddata <= 8'h53;
            13'h0398: rddata <= 8'h54;
            13'h0399: rddata <= 8'h43;
            13'h039A: rddata <= 8'h4E;
            13'h039B: rddata <= 8'h55;
            13'h039C: rddata <= 8'h46;
            13'h039D: rddata <= 8'h4D;
            13'h039E: rddata <= 8'h4F;
            13'h039F: rddata <= 8'h21;
            13'h03A0: rddata <= 8'h04;
            13'h03A1: rddata <= 8'h00;
            13'h03A2: rddata <= 8'h39;
            13'h03A3: rddata <= 8'h7E;
            13'h03A4: rddata <= 8'h23;
            13'h03A5: rddata <= 8'hFE;
            13'h03A6: rddata <= 8'h81;
            13'h03A7: rddata <= 8'hC0;
            13'h03A8: rddata <= 8'h4E;
            13'h03A9: rddata <= 8'h23;
            13'h03AA: rddata <= 8'h46;
            13'h03AB: rddata <= 8'h23;
            13'h03AC: rddata <= 8'hE5;
            13'h03AD: rddata <= 8'h60;
            13'h03AE: rddata <= 8'h69;
            13'h03AF: rddata <= 8'h7A;
            13'h03B0: rddata <= 8'hB3;
            13'h03B1: rddata <= 8'hEB;
            13'h03B2: rddata <= 8'h28;
            13'h03B3: rddata <= 8'h02;
            13'h03B4: rddata <= 8'hEB;
            13'h03B5: rddata <= 8'hE7;
            13'h03B6: rddata <= 8'h01;
            13'h03B7: rddata <= 8'h0D;
            13'h03B8: rddata <= 8'h00;
            13'h03B9: rddata <= 8'hE1;
            13'h03BA: rddata <= 8'hC8;
            13'h03BB: rddata <= 8'h09;
            13'h03BC: rddata <= 8'h18;
            13'h03BD: rddata <= 8'hE5;
            13'h03BE: rddata <= 8'h2A;
            13'h03BF: rddata <= 8'hC9;
            13'h03C0: rddata <= 8'h38;
            13'h03C1: rddata <= 8'h22;
            13'h03C2: rddata <= 8'h4D;
            13'h03C3: rddata <= 8'h38;
            13'h03C4: rddata <= 8'h1E;
            13'h03C5: rddata <= 8'h02;
            13'h03C6: rddata <= 8'h01;
            13'h03C7: rddata <= 8'h1E;
            13'h03C8: rddata <= 8'h14;
            13'h03C9: rddata <= 8'h01;
            13'h03CA: rddata <= 8'h1E;
            13'h03CB: rddata <= 8'h00;
            13'h03CC: rddata <= 8'h01;
            13'h03CD: rddata <= 8'h1E;
            13'h03CE: rddata <= 8'h12;
            13'h03CF: rddata <= 8'h01;
            13'h03D0: rddata <= 8'h1E;
            13'h03D1: rddata <= 8'h22;
            13'h03D2: rddata <= 8'h01;
            13'h03D3: rddata <= 8'h1E;
            13'h03D4: rddata <= 8'h0A;
            13'h03D5: rddata <= 8'h01;
            13'h03D6: rddata <= 8'h1E;
            13'h03D7: rddata <= 8'h24;
            13'h03D8: rddata <= 8'h01;
            13'h03D9: rddata <= 8'h1E;
            13'h03DA: rddata <= 8'h18;
            13'h03DB: rddata <= 8'hCD;
            13'h03DC: rddata <= 8'hE5;
            13'h03DD: rddata <= 8'h0B;
            13'h03DE: rddata <= 8'hF7;
            13'h03DF: rddata <= 8'h00;
            13'h03E0: rddata <= 8'hCD;
            13'h03E1: rddata <= 8'hDE;
            13'h03E2: rddata <= 8'h19;
            13'h03E3: rddata <= 8'h21;
            13'h03E4: rddata <= 8'h79;
            13'h03E5: rddata <= 8'h03;
            13'h03E6: rddata <= 8'hF7;
            13'h03E7: rddata <= 8'h01;
            13'h03E8: rddata <= 8'h57;
            13'h03E9: rddata <= 8'h19;
            13'h03EA: rddata <= 8'h3E;
            13'h03EB: rddata <= 8'h3F;
            13'h03EC: rddata <= 8'hDF;
            13'h03ED: rddata <= 8'h7E;
            13'h03EE: rddata <= 8'hDF;
            13'h03EF: rddata <= 8'hD7;
            13'h03F0: rddata <= 8'hDF;
            13'h03F1: rddata <= 8'h21;
            13'h03F2: rddata <= 8'h61;
            13'h03F3: rddata <= 8'h03;
            13'h03F4: rddata <= 8'hCD;
            13'h03F5: rddata <= 8'h9D;
            13'h03F6: rddata <= 8'h0E;
            13'h03F7: rddata <= 8'h2A;
            13'h03F8: rddata <= 8'h4D;
            13'h03F9: rddata <= 8'h38;
            13'h03FA: rddata <= 8'h7C;
            13'h03FB: rddata <= 8'hA5;
            13'h03FC: rddata <= 8'h3C;
            13'h03FD: rddata <= 8'hC4;
            13'h03FE: rddata <= 8'h6D;
            13'h03FF: rddata <= 8'h16;
            13'h0400: rddata <= 8'h3E;
            13'h0401: rddata <= 8'hC1;
            13'h0402: rddata <= 8'hF7;
            13'h0403: rddata <= 8'h02;
            13'h0404: rddata <= 8'hCD;
            13'h0405: rddata <= 8'hBE;
            13'h0406: rddata <= 8'h19;
            13'h0407: rddata <= 8'hAF;
            13'h0408: rddata <= 8'h32;
            13'h0409: rddata <= 8'h08;
            13'h040A: rddata <= 8'h38;
            13'h040B: rddata <= 8'hCD;
            13'h040C: rddata <= 8'hDE;
            13'h040D: rddata <= 8'h19;
            13'h040E: rddata <= 8'h21;
            13'h040F: rddata <= 8'h6E;
            13'h0410: rddata <= 8'h03;
            13'h0411: rddata <= 8'hCD;
            13'h0412: rddata <= 8'h9D;
            13'h0413: rddata <= 8'h0E;
            13'h0414: rddata <= 8'h21;
            13'h0415: rddata <= 8'hFF;
            13'h0416: rddata <= 8'hFF;
            13'h0417: rddata <= 8'h22;
            13'h0418: rddata <= 8'h4D;
            13'h0419: rddata <= 8'h38;
            13'h041A: rddata <= 8'hCD;
            13'h041B: rddata <= 8'h85;
            13'h041C: rddata <= 8'h0D;
            13'h041D: rddata <= 8'h38;
            13'h041E: rddata <= 8'hF5;
            13'h041F: rddata <= 8'hD7;
            13'h0420: rddata <= 8'h3C;
            13'h0421: rddata <= 8'h3D;
            13'h0422: rddata <= 8'h28;
            13'h0423: rddata <= 8'hF0;
            13'h0424: rddata <= 8'hF5;
            13'h0425: rddata <= 8'hCD;
            13'h0426: rddata <= 8'h9C;
            13'h0427: rddata <= 8'h06;
            13'h0428: rddata <= 8'hD5;
            13'h0429: rddata <= 8'hCD;
            13'h042A: rddata <= 8'hBC;
            13'h042B: rddata <= 8'h04;
            13'h042C: rddata <= 8'h47;
            13'h042D: rddata <= 8'hD1;
            13'h042E: rddata <= 8'hF1;
            13'h042F: rddata <= 8'hF7;
            13'h0430: rddata <= 8'h03;
            13'h0431: rddata <= 8'hD2;
            13'h0432: rddata <= 8'h4B;
            13'h0433: rddata <= 8'h06;
            13'h0434: rddata <= 8'hD5;
            13'h0435: rddata <= 8'hC5;
            13'h0436: rddata <= 8'hAF;
            13'h0437: rddata <= 8'h32;
            13'h0438: rddata <= 8'hCC;
            13'h0439: rddata <= 8'h38;
            13'h043A: rddata <= 8'hD7;
            13'h043B: rddata <= 8'hB7;
            13'h043C: rddata <= 8'hF5;
            13'h043D: rddata <= 8'hCD;
            13'h043E: rddata <= 8'h9F;
            13'h043F: rddata <= 8'h04;
            13'h0440: rddata <= 8'h38;
            13'h0441: rddata <= 8'h06;
            13'h0442: rddata <= 8'hF1;
            13'h0443: rddata <= 8'hF5;
            13'h0444: rddata <= 8'hCA;
            13'h0445: rddata <= 8'hF3;
            13'h0446: rddata <= 8'h06;
            13'h0447: rddata <= 8'hB7;
            13'h0448: rddata <= 8'hC5;
            13'h0449: rddata <= 8'h30;
            13'h044A: rddata <= 8'h10;
            13'h044B: rddata <= 8'hEB;
            13'h044C: rddata <= 8'h2A;
            13'h044D: rddata <= 8'hD6;
            13'h044E: rddata <= 8'h38;
            13'h044F: rddata <= 8'h1A;
            13'h0450: rddata <= 8'h02;
            13'h0451: rddata <= 8'h03;
            13'h0452: rddata <= 8'h13;
            13'h0453: rddata <= 8'hE7;
            13'h0454: rddata <= 8'h20;
            13'h0455: rddata <= 8'hF9;
            13'h0456: rddata <= 8'h60;
            13'h0457: rddata <= 8'h69;
            13'h0458: rddata <= 8'h22;
            13'h0459: rddata <= 8'hD6;
            13'h045A: rddata <= 8'h38;
            13'h045B: rddata <= 8'hD1;
            13'h045C: rddata <= 8'hF1;
            13'h045D: rddata <= 8'h28;
            13'h045E: rddata <= 8'h21;
            13'h045F: rddata <= 8'h2A;
            13'h0460: rddata <= 8'hD6;
            13'h0461: rddata <= 8'h38;
            13'h0462: rddata <= 8'hE3;
            13'h0463: rddata <= 8'hC1;
            13'h0464: rddata <= 8'h09;
            13'h0465: rddata <= 8'hE5;
            13'h0466: rddata <= 8'hCD;
            13'h0467: rddata <= 8'h92;
            13'h0468: rddata <= 8'h0B;
            13'h0469: rddata <= 8'hE1;
            13'h046A: rddata <= 8'h22;
            13'h046B: rddata <= 8'hD6;
            13'h046C: rddata <= 8'h38;
            13'h046D: rddata <= 8'hEB;
            13'h046E: rddata <= 8'h74;
            13'h046F: rddata <= 8'hD1;
            13'h0470: rddata <= 8'h23;
            13'h0471: rddata <= 8'h23;
            13'h0472: rddata <= 8'h73;
            13'h0473: rddata <= 8'h23;
            13'h0474: rddata <= 8'h72;
            13'h0475: rddata <= 8'h23;
            13'h0476: rddata <= 8'h11;
            13'h0477: rddata <= 8'h60;
            13'h0478: rddata <= 8'h38;
            13'h0479: rddata <= 8'h1A;
            13'h047A: rddata <= 8'h77;
            13'h047B: rddata <= 8'h23;
            13'h047C: rddata <= 8'h13;
            13'h047D: rddata <= 8'hB7;
            13'h047E: rddata <= 8'h20;
            13'h047F: rddata <= 8'hF9;
            13'h0480: rddata <= 8'hF7;
            13'h0481: rddata <= 8'h04;
            13'h0482: rddata <= 8'hCD;
            13'h0483: rddata <= 8'hCB;
            13'h0484: rddata <= 8'h0B;
            13'h0485: rddata <= 8'hF7;
            13'h0486: rddata <= 8'h05;
            13'h0487: rddata <= 8'h23;
            13'h0488: rddata <= 8'hEB;
            13'h0489: rddata <= 8'h62;
            13'h048A: rddata <= 8'h6B;
            13'h048B: rddata <= 8'h7E;
            13'h048C: rddata <= 8'h23;
            13'h048D: rddata <= 8'hB6;
            13'h048E: rddata <= 8'hCA;
            13'h048F: rddata <= 8'h14;
            13'h0490: rddata <= 8'h04;
            13'h0491: rddata <= 8'h23;
            13'h0492: rddata <= 8'h23;
            13'h0493: rddata <= 8'h23;
            13'h0494: rddata <= 8'hAF;
            13'h0495: rddata <= 8'hBE;
            13'h0496: rddata <= 8'h23;
            13'h0497: rddata <= 8'h20;
            13'h0498: rddata <= 8'hFC;
            13'h0499: rddata <= 8'hEB;
            13'h049A: rddata <= 8'h73;
            13'h049B: rddata <= 8'h23;
            13'h049C: rddata <= 8'h72;
            13'h049D: rddata <= 8'h18;
            13'h049E: rddata <= 8'hEA;
            13'h049F: rddata <= 8'h2A;
            13'h04A0: rddata <= 8'h4F;
            13'h04A1: rddata <= 8'h38;
            13'h04A2: rddata <= 8'h44;
            13'h04A3: rddata <= 8'h4D;
            13'h04A4: rddata <= 8'h7E;
            13'h04A5: rddata <= 8'h23;
            13'h04A6: rddata <= 8'hB6;
            13'h04A7: rddata <= 8'h2B;
            13'h04A8: rddata <= 8'hC8;
            13'h04A9: rddata <= 8'h23;
            13'h04AA: rddata <= 8'h23;
            13'h04AB: rddata <= 8'h7E;
            13'h04AC: rddata <= 8'h23;
            13'h04AD: rddata <= 8'h66;
            13'h04AE: rddata <= 8'h6F;
            13'h04AF: rddata <= 8'hE7;
            13'h04B0: rddata <= 8'h60;
            13'h04B1: rddata <= 8'h69;
            13'h04B2: rddata <= 8'h7E;
            13'h04B3: rddata <= 8'h23;
            13'h04B4: rddata <= 8'h66;
            13'h04B5: rddata <= 8'h6F;
            13'h04B6: rddata <= 8'h3F;
            13'h04B7: rddata <= 8'hC8;
            13'h04B8: rddata <= 8'h3F;
            13'h04B9: rddata <= 8'hD0;
            13'h04BA: rddata <= 8'h18;
            13'h04BB: rddata <= 8'hE6;
            13'h04BC: rddata <= 8'hAF;
            13'h04BD: rddata <= 8'h32;
            13'h04BE: rddata <= 8'hAC;
            13'h04BF: rddata <= 8'h38;
            13'h04C0: rddata <= 8'h0E;
            13'h04C1: rddata <= 8'h05;
            13'h04C2: rddata <= 8'h11;
            13'h04C3: rddata <= 8'h60;
            13'h04C4: rddata <= 8'h38;
            13'h04C5: rddata <= 8'h7E;
            13'h04C6: rddata <= 8'hFE;
            13'h04C7: rddata <= 8'h20;
            13'h04C8: rddata <= 8'hCA;
            13'h04C9: rddata <= 8'h3C;
            13'h04CA: rddata <= 8'h05;
            13'h04CB: rddata <= 8'h47;
            13'h04CC: rddata <= 8'hFE;
            13'h04CD: rddata <= 8'h22;
            13'h04CE: rddata <= 8'hCA;
            13'h04CF: rddata <= 8'h58;
            13'h04D0: rddata <= 8'h05;
            13'h04D1: rddata <= 8'hB7;
            13'h04D2: rddata <= 8'hCA;
            13'h04D3: rddata <= 8'h5E;
            13'h04D4: rddata <= 8'h05;
            13'h04D5: rddata <= 8'h3A;
            13'h04D6: rddata <= 8'hAC;
            13'h04D7: rddata <= 8'h38;
            13'h04D8: rddata <= 8'hB7;
            13'h04D9: rddata <= 8'h7E;
            13'h04DA: rddata <= 8'hC2;
            13'h04DB: rddata <= 8'h3C;
            13'h04DC: rddata <= 8'h05;
            13'h04DD: rddata <= 8'hFE;
            13'h04DE: rddata <= 8'h3F;
            13'h04DF: rddata <= 8'h3E;
            13'h04E0: rddata <= 8'h95;
            13'h04E1: rddata <= 8'hCA;
            13'h04E2: rddata <= 8'h3C;
            13'h04E3: rddata <= 8'h05;
            13'h04E4: rddata <= 8'h7E;
            13'h04E5: rddata <= 8'hFE;
            13'h04E6: rddata <= 8'h30;
            13'h04E7: rddata <= 8'h38;
            13'h04E8: rddata <= 8'h05;
            13'h04E9: rddata <= 8'hFE;
            13'h04EA: rddata <= 8'h3C;
            13'h04EB: rddata <= 8'hDA;
            13'h04EC: rddata <= 8'h3C;
            13'h04ED: rddata <= 8'h05;
            13'h04EE: rddata <= 8'hD5;
            13'h04EF: rddata <= 8'h11;
            13'h04F0: rddata <= 8'h44;
            13'h04F1: rddata <= 8'h02;
            13'h04F2: rddata <= 8'hC5;
            13'h04F3: rddata <= 8'h01;
            13'h04F4: rddata <= 8'h36;
            13'h04F5: rddata <= 8'h05;
            13'h04F6: rddata <= 8'hC5;
            13'h04F7: rddata <= 8'h06;
            13'h04F8: rddata <= 8'h7F;
            13'h04F9: rddata <= 8'h7E;
            13'h04FA: rddata <= 8'hFE;
            13'h04FB: rddata <= 8'h61;
            13'h04FC: rddata <= 8'h38;
            13'h04FD: rddata <= 8'h07;
            13'h04FE: rddata <= 8'hFE;
            13'h04FF: rddata <= 8'h7B;
            13'h0500: rddata <= 8'h30;
            13'h0501: rddata <= 8'h03;
            13'h0502: rddata <= 8'hE6;
            13'h0503: rddata <= 8'h5F;
            13'h0504: rddata <= 8'h77;
            13'h0505: rddata <= 8'h4E;
            13'h0506: rddata <= 8'hEB;
            13'h0507: rddata <= 8'h23;
            13'h0508: rddata <= 8'hB6;
            13'h0509: rddata <= 8'hF2;
            13'h050A: rddata <= 8'h07;
            13'h050B: rddata <= 8'h05;
            13'h050C: rddata <= 8'h04;
            13'h050D: rddata <= 8'h7E;
            13'h050E: rddata <= 8'hE6;
            13'h050F: rddata <= 8'h7F;
            13'h0510: rddata <= 8'hC8;
            13'h0511: rddata <= 8'hB9;
            13'h0512: rddata <= 8'h20;
            13'h0513: rddata <= 8'hF3;
            13'h0514: rddata <= 8'hEB;
            13'h0515: rddata <= 8'hE5;
            13'h0516: rddata <= 8'h13;
            13'h0517: rddata <= 8'h1A;
            13'h0518: rddata <= 8'hB7;
            13'h0519: rddata <= 8'hFA;
            13'h051A: rddata <= 8'h32;
            13'h051B: rddata <= 8'h05;
            13'h051C: rddata <= 8'h4F;
            13'h051D: rddata <= 8'h78;
            13'h051E: rddata <= 8'hFE;
            13'h051F: rddata <= 8'h88;
            13'h0520: rddata <= 8'h20;
            13'h0521: rddata <= 8'h02;
            13'h0522: rddata <= 8'hD7;
            13'h0523: rddata <= 8'h2B;
            13'h0524: rddata <= 8'h23;
            13'h0525: rddata <= 8'h7E;
            13'h0526: rddata <= 8'hFE;
            13'h0527: rddata <= 8'h61;
            13'h0528: rddata <= 8'h38;
            13'h0529: rddata <= 8'h02;
            13'h052A: rddata <= 8'hE6;
            13'h052B: rddata <= 8'h5F;
            13'h052C: rddata <= 8'hB9;
            13'h052D: rddata <= 8'h28;
            13'h052E: rddata <= 8'hE7;
            13'h052F: rddata <= 8'hE1;
            13'h0530: rddata <= 8'h18;
            13'h0531: rddata <= 8'hD3;
            13'h0532: rddata <= 8'h48;
            13'h0533: rddata <= 8'hF1;
            13'h0534: rddata <= 8'hEB;
            13'h0535: rddata <= 8'hC9;
            13'h0536: rddata <= 8'hF7;
            13'h0537: rddata <= 8'h0A;
            13'h0538: rddata <= 8'hEB;
            13'h0539: rddata <= 8'h79;
            13'h053A: rddata <= 8'hC1;
            13'h053B: rddata <= 8'hD1;
            13'h053C: rddata <= 8'h23;
            13'h053D: rddata <= 8'h12;
            13'h053E: rddata <= 8'h13;
            13'h053F: rddata <= 8'h0C;
            13'h0540: rddata <= 8'hD6;
            13'h0541: rddata <= 8'h3A;
            13'h0542: rddata <= 8'h28;
            13'h0543: rddata <= 8'h04;
            13'h0544: rddata <= 8'hFE;
            13'h0545: rddata <= 8'h49;
            13'h0546: rddata <= 8'h20;
            13'h0547: rddata <= 8'h03;
            13'h0548: rddata <= 8'h32;
            13'h0549: rddata <= 8'hAC;
            13'h054A: rddata <= 8'h38;
            13'h054B: rddata <= 8'hD6;
            13'h054C: rddata <= 8'h54;
            13'h054D: rddata <= 8'hC2;
            13'h054E: rddata <= 8'hC5;
            13'h054F: rddata <= 8'h04;
            13'h0550: rddata <= 8'h47;
            13'h0551: rddata <= 8'h7E;
            13'h0552: rddata <= 8'hB7;
            13'h0553: rddata <= 8'h28;
            13'h0554: rddata <= 8'h09;
            13'h0555: rddata <= 8'hB8;
            13'h0556: rddata <= 8'h28;
            13'h0557: rddata <= 8'hE4;
            13'h0558: rddata <= 8'h23;
            13'h0559: rddata <= 8'h12;
            13'h055A: rddata <= 8'h0C;
            13'h055B: rddata <= 8'h13;
            13'h055C: rddata <= 8'h18;
            13'h055D: rddata <= 8'hF3;
            13'h055E: rddata <= 8'h21;
            13'h055F: rddata <= 8'h5F;
            13'h0560: rddata <= 8'h38;
            13'h0561: rddata <= 8'h12;
            13'h0562: rddata <= 8'h13;
            13'h0563: rddata <= 8'h12;
            13'h0564: rddata <= 8'h13;
            13'h0565: rddata <= 8'h12;
            13'h0566: rddata <= 8'hC9;
            13'h0567: rddata <= 8'h3E;
            13'h0568: rddata <= 8'h01;
            13'h0569: rddata <= 8'h32;
            13'h056A: rddata <= 8'h47;
            13'h056B: rddata <= 8'h38;
            13'h056C: rddata <= 8'h3E;
            13'h056D: rddata <= 8'h17;
            13'h056E: rddata <= 8'h32;
            13'h056F: rddata <= 8'h08;
            13'h0570: rddata <= 8'h38;
            13'h0571: rddata <= 8'hCD;
            13'h0572: rddata <= 8'h9C;
            13'h0573: rddata <= 8'h06;
            13'h0574: rddata <= 8'hC0;
            13'h0575: rddata <= 8'hC1;
            13'h0576: rddata <= 8'hCD;
            13'h0577: rddata <= 8'h9F;
            13'h0578: rddata <= 8'h04;
            13'h0579: rddata <= 8'hC5;
            13'h057A: rddata <= 8'hE1;
            13'h057B: rddata <= 8'h4E;
            13'h057C: rddata <= 8'h23;
            13'h057D: rddata <= 8'h46;
            13'h057E: rddata <= 8'h23;
            13'h057F: rddata <= 8'h78;
            13'h0580: rddata <= 8'hB1;
            13'h0581: rddata <= 8'hCA;
            13'h0582: rddata <= 8'h02;
            13'h0583: rddata <= 8'h04;
            13'h0584: rddata <= 8'hCD;
            13'h0585: rddata <= 8'h25;
            13'h0586: rddata <= 8'h1A;
            13'h0587: rddata <= 8'hC5;
            13'h0588: rddata <= 8'hCD;
            13'h0589: rddata <= 8'hEA;
            13'h058A: rddata <= 8'h19;
            13'h058B: rddata <= 8'h5E;
            13'h058C: rddata <= 8'h23;
            13'h058D: rddata <= 8'h56;
            13'h058E: rddata <= 8'h23;
            13'h058F: rddata <= 8'hE5;
            13'h0590: rddata <= 8'hEB;
            13'h0591: rddata <= 8'hCD;
            13'h0592: rddata <= 8'h75;
            13'h0593: rddata <= 8'h16;
            13'h0594: rddata <= 8'h3E;
            13'h0595: rddata <= 8'h20;
            13'h0596: rddata <= 8'hE1;
            13'h0597: rddata <= 8'hDF;
            13'h0598: rddata <= 8'h7E;
            13'h0599: rddata <= 8'h23;
            13'h059A: rddata <= 8'hB7;
            13'h059B: rddata <= 8'h28;
            13'h059C: rddata <= 8'hDD;
            13'h059D: rddata <= 8'hF2;
            13'h059E: rddata <= 8'h97;
            13'h059F: rddata <= 8'h05;
            13'h05A0: rddata <= 8'hF7;
            13'h05A1: rddata <= 8'h16;
            13'h05A2: rddata <= 8'hD6;
            13'h05A3: rddata <= 8'h7F;
            13'h05A4: rddata <= 8'h4F;
            13'h05A5: rddata <= 8'h11;
            13'h05A6: rddata <= 8'h45;
            13'h05A7: rddata <= 8'h02;
            13'h05A8: rddata <= 8'h1A;
            13'h05A9: rddata <= 8'h13;
            13'h05AA: rddata <= 8'hB7;
            13'h05AB: rddata <= 8'hF2;
            13'h05AC: rddata <= 8'hA8;
            13'h05AD: rddata <= 8'h05;
            13'h05AE: rddata <= 8'h0D;
            13'h05AF: rddata <= 8'h20;
            13'h05B0: rddata <= 8'hF7;
            13'h05B1: rddata <= 8'hE6;
            13'h05B2: rddata <= 8'h7F;
            13'h05B3: rddata <= 8'hDF;
            13'h05B4: rddata <= 8'h1A;
            13'h05B5: rddata <= 8'h13;
            13'h05B6: rddata <= 8'hB7;
            13'h05B7: rddata <= 8'hF2;
            13'h05B8: rddata <= 8'hB1;
            13'h05B9: rddata <= 8'h05;
            13'h05BA: rddata <= 8'h18;
            13'h05BB: rddata <= 8'hDC;
            13'h05BC: rddata <= 8'h3E;
            13'h05BD: rddata <= 8'h64;
            13'h05BE: rddata <= 8'h32;
            13'h05BF: rddata <= 8'hCB;
            13'h05C0: rddata <= 8'h38;
            13'h05C1: rddata <= 8'hCD;
            13'h05C2: rddata <= 8'h31;
            13'h05C3: rddata <= 8'h07;
            13'h05C4: rddata <= 8'hC1;
            13'h05C5: rddata <= 8'hE5;
            13'h05C6: rddata <= 8'hCD;
            13'h05C7: rddata <= 8'h1C;
            13'h05C8: rddata <= 8'h07;
            13'h05C9: rddata <= 8'h22;
            13'h05CA: rddata <= 8'hC7;
            13'h05CB: rddata <= 8'h38;
            13'h05CC: rddata <= 8'h21;
            13'h05CD: rddata <= 8'h02;
            13'h05CE: rddata <= 8'h00;
            13'h05CF: rddata <= 8'h39;
            13'h05D0: rddata <= 8'hCD;
            13'h05D1: rddata <= 8'hA3;
            13'h05D2: rddata <= 8'h03;
            13'h05D3: rddata <= 8'h20;
            13'h05D4: rddata <= 8'h14;
            13'h05D5: rddata <= 8'h09;
            13'h05D6: rddata <= 8'hD5;
            13'h05D7: rddata <= 8'h2B;
            13'h05D8: rddata <= 8'h56;
            13'h05D9: rddata <= 8'h2B;
            13'h05DA: rddata <= 8'h5E;
            13'h05DB: rddata <= 8'h23;
            13'h05DC: rddata <= 8'h23;
            13'h05DD: rddata <= 8'hE5;
            13'h05DE: rddata <= 8'h2A;
            13'h05DF: rddata <= 8'hC7;
            13'h05E0: rddata <= 8'h38;
            13'h05E1: rddata <= 8'hE7;
            13'h05E2: rddata <= 8'hE1;
            13'h05E3: rddata <= 8'hD1;
            13'h05E4: rddata <= 8'h20;
            13'h05E5: rddata <= 8'hEA;
            13'h05E6: rddata <= 8'hD1;
            13'h05E7: rddata <= 8'hF9;
            13'h05E8: rddata <= 8'h0C;
            13'h05E9: rddata <= 8'hD1;
            13'h05EA: rddata <= 8'hEB;
            13'h05EB: rddata <= 8'h0E;
            13'h05EC: rddata <= 8'h08;
            13'h05ED: rddata <= 8'hCD;
            13'h05EE: rddata <= 8'hA0;
            13'h05EF: rddata <= 8'h0B;
            13'h05F0: rddata <= 8'hE5;
            13'h05F1: rddata <= 8'h2A;
            13'h05F2: rddata <= 8'hC7;
            13'h05F3: rddata <= 8'h38;
            13'h05F4: rddata <= 8'hE3;
            13'h05F5: rddata <= 8'hE5;
            13'h05F6: rddata <= 8'h2A;
            13'h05F7: rddata <= 8'h4D;
            13'h05F8: rddata <= 8'h38;
            13'h05F9: rddata <= 8'hE3;
            13'h05FA: rddata <= 8'hCD;
            13'h05FB: rddata <= 8'h75;
            13'h05FC: rddata <= 8'h09;
            13'h05FD: rddata <= 8'hCF;
            13'h05FE: rddata <= 8'hA1;
            13'h05FF: rddata <= 8'hCD;
            13'h0600: rddata <= 8'h72;
            13'h0601: rddata <= 8'h09;
            13'h0602: rddata <= 8'hE5;
            13'h0603: rddata <= 8'hCD;
            13'h0604: rddata <= 8'h2E;
            13'h0605: rddata <= 8'h15;
            13'h0606: rddata <= 8'hE1;
            13'h0607: rddata <= 8'hC5;
            13'h0608: rddata <= 8'hD5;
            13'h0609: rddata <= 8'h01;
            13'h060A: rddata <= 8'h00;
            13'h060B: rddata <= 8'h81;
            13'h060C: rddata <= 8'h51;
            13'h060D: rddata <= 8'h5A;
            13'h060E: rddata <= 8'h7E;
            13'h060F: rddata <= 8'hFE;
            13'h0610: rddata <= 8'hA7;
            13'h0611: rddata <= 8'h3E;
            13'h0612: rddata <= 8'h01;
            13'h0613: rddata <= 8'h20;
            13'h0614: rddata <= 8'h0A;
            13'h0615: rddata <= 8'hD7;
            13'h0616: rddata <= 8'hCD;
            13'h0617: rddata <= 8'h72;
            13'h0618: rddata <= 8'h09;
            13'h0619: rddata <= 8'hE5;
            13'h061A: rddata <= 8'hCD;
            13'h061B: rddata <= 8'h2E;
            13'h061C: rddata <= 8'h15;
            13'h061D: rddata <= 8'hEF;
            13'h061E: rddata <= 8'hE1;
            13'h061F: rddata <= 8'hC5;
            13'h0620: rddata <= 8'hD5;
            13'h0621: rddata <= 8'hF5;
            13'h0622: rddata <= 8'h33;
            13'h0623: rddata <= 8'hE5;
            13'h0624: rddata <= 8'h2A;
            13'h0625: rddata <= 8'hCE;
            13'h0626: rddata <= 8'h38;
            13'h0627: rddata <= 8'hE3;
            13'h0628: rddata <= 8'h06;
            13'h0629: rddata <= 8'h81;
            13'h062A: rddata <= 8'hC5;
            13'h062B: rddata <= 8'h33;
            13'h062C: rddata <= 8'h22;
            13'h062D: rddata <= 8'hCE;
            13'h062E: rddata <= 8'h38;
            13'h062F: rddata <= 8'hCD;
            13'h0630: rddata <= 8'hC2;
            13'h0631: rddata <= 8'h1F;
            13'h0632: rddata <= 8'h7E;
            13'h0633: rddata <= 8'hFE;
            13'h0634: rddata <= 8'h3A;
            13'h0635: rddata <= 8'h28;
            13'h0636: rddata <= 8'h14;
            13'h0637: rddata <= 8'hB7;
            13'h0638: rddata <= 8'hC2;
            13'h0639: rddata <= 8'hC4;
            13'h063A: rddata <= 8'h03;
            13'h063B: rddata <= 8'h23;
            13'h063C: rddata <= 8'h7E;
            13'h063D: rddata <= 8'h23;
            13'h063E: rddata <= 8'hB6;
            13'h063F: rddata <= 8'hCA;
            13'h0640: rddata <= 8'h29;
            13'h0641: rddata <= 8'h0C;
            13'h0642: rddata <= 8'h23;
            13'h0643: rddata <= 8'h5E;
            13'h0644: rddata <= 8'h23;
            13'h0645: rddata <= 8'h56;
            13'h0646: rddata <= 8'hEB;
            13'h0647: rddata <= 8'h22;
            13'h0648: rddata <= 8'h4D;
            13'h0649: rddata <= 8'h38;
            13'h064A: rddata <= 8'hEB;
            13'h064B: rddata <= 8'hD7;
            13'h064C: rddata <= 8'h11;
            13'h064D: rddata <= 8'h2C;
            13'h064E: rddata <= 8'h06;
            13'h064F: rddata <= 8'hD5;
            13'h0650: rddata <= 8'hC8;
            13'h0651: rddata <= 8'hD6;
            13'h0652: rddata <= 8'h80;
            13'h0653: rddata <= 8'hDA;
            13'h0654: rddata <= 8'h31;
            13'h0655: rddata <= 8'h07;
            13'h0656: rddata <= 8'hFE;
            13'h0657: rddata <= 8'h20;
            13'h0658: rddata <= 8'hF7;
            13'h0659: rddata <= 8'h17;
            13'h065A: rddata <= 8'hD2;
            13'h065B: rddata <= 8'hC4;
            13'h065C: rddata <= 8'h03;
            13'h065D: rddata <= 8'h07;
            13'h065E: rddata <= 8'h4F;
            13'h065F: rddata <= 8'h06;
            13'h0660: rddata <= 8'h00;
            13'h0661: rddata <= 8'hEB;
            13'h0662: rddata <= 8'h21;
            13'h0663: rddata <= 8'hD5;
            13'h0664: rddata <= 8'h01;
            13'h0665: rddata <= 8'h09;
            13'h0666: rddata <= 8'h4E;
            13'h0667: rddata <= 8'h23;
            13'h0668: rddata <= 8'h46;
            13'h0669: rddata <= 8'hC5;
            13'h066A: rddata <= 8'hEB;
            13'h066B: rddata <= 8'h23;
            13'h066C: rddata <= 8'h7E;
            13'h066D: rddata <= 8'hFE;
            13'h066E: rddata <= 8'h3A;
            13'h066F: rddata <= 8'hD0;
            13'h0670: rddata <= 8'hFE;
            13'h0671: rddata <= 8'h20;
            13'h0672: rddata <= 8'h28;
            13'h0673: rddata <= 8'hF7;
            13'h0674: rddata <= 8'hFE;
            13'h0675: rddata <= 8'h30;
            13'h0676: rddata <= 8'h3F;
            13'h0677: rddata <= 8'h3C;
            13'h0678: rddata <= 8'h3D;
            13'h0679: rddata <= 8'hC9;
            13'h067A: rddata <= 8'hD7;
            13'h067B: rddata <= 8'hCD;
            13'h067C: rddata <= 8'h72;
            13'h067D: rddata <= 8'h09;
            13'h067E: rddata <= 8'hEF;
            13'h067F: rddata <= 8'hFA;
            13'h0680: rddata <= 8'h97;
            13'h0681: rddata <= 8'h06;
            13'h0682: rddata <= 8'h3A;
            13'h0683: rddata <= 8'hE7;
            13'h0684: rddata <= 8'h38;
            13'h0685: rddata <= 8'hFE;
            13'h0686: rddata <= 8'h90;
            13'h0687: rddata <= 8'hDA;
            13'h0688: rddata <= 8'h86;
            13'h0689: rddata <= 8'h15;
            13'h068A: rddata <= 8'h01;
            13'h068B: rddata <= 8'h80;
            13'h068C: rddata <= 8'h90;
            13'h068D: rddata <= 8'h11;
            13'h068E: rddata <= 8'h00;
            13'h068F: rddata <= 8'h00;
            13'h0690: rddata <= 8'hE5;
            13'h0691: rddata <= 8'hCD;
            13'h0692: rddata <= 8'h5B;
            13'h0693: rddata <= 8'h15;
            13'h0694: rddata <= 8'hE1;
            13'h0695: rddata <= 8'h51;
            13'h0696: rddata <= 8'hC8;
            13'h0697: rddata <= 8'h1E;
            13'h0698: rddata <= 8'h08;
            13'h0699: rddata <= 8'hC3;
            13'h069A: rddata <= 8'hDB;
            13'h069B: rddata <= 8'h03;
            13'h069C: rddata <= 8'h2B;
            13'h069D: rddata <= 8'h11;
            13'h069E: rddata <= 8'h00;
            13'h069F: rddata <= 8'h00;
            13'h06A0: rddata <= 8'hD7;
            13'h06A1: rddata <= 8'hD0;
            13'h06A2: rddata <= 8'hE5;
            13'h06A3: rddata <= 8'hF5;
            13'h06A4: rddata <= 8'h21;
            13'h06A5: rddata <= 8'h98;
            13'h06A6: rddata <= 8'h19;
            13'h06A7: rddata <= 8'hE7;
            13'h06A8: rddata <= 8'h38;
            13'h06A9: rddata <= 8'h11;
            13'h06AA: rddata <= 8'h62;
            13'h06AB: rddata <= 8'h6B;
            13'h06AC: rddata <= 8'h19;
            13'h06AD: rddata <= 8'h29;
            13'h06AE: rddata <= 8'h19;
            13'h06AF: rddata <= 8'h29;
            13'h06B0: rddata <= 8'hF1;
            13'h06B1: rddata <= 8'hD6;
            13'h06B2: rddata <= 8'h30;
            13'h06B3: rddata <= 8'h5F;
            13'h06B4: rddata <= 8'h16;
            13'h06B5: rddata <= 8'h00;
            13'h06B6: rddata <= 8'h19;
            13'h06B7: rddata <= 8'hEB;
            13'h06B8: rddata <= 8'hE1;
            13'h06B9: rddata <= 8'h18;
            13'h06BA: rddata <= 8'hE5;
            13'h06BB: rddata <= 8'hF1;
            13'h06BC: rddata <= 8'hE1;
            13'h06BD: rddata <= 8'hC9;
            13'h06BE: rddata <= 8'hF7;
            13'h06BF: rddata <= 8'h18;
            13'h06C0: rddata <= 8'hCA;
            13'h06C1: rddata <= 8'hCB;
            13'h06C2: rddata <= 8'h0B;
            13'h06C3: rddata <= 8'hCD;
            13'h06C4: rddata <= 8'hCF;
            13'h06C5: rddata <= 8'h0B;
            13'h06C6: rddata <= 8'h01;
            13'h06C7: rddata <= 8'h2C;
            13'h06C8: rddata <= 8'h06;
            13'h06C9: rddata <= 8'h18;
            13'h06CA: rddata <= 8'h10;
            13'h06CB: rddata <= 8'h0E;
            13'h06CC: rddata <= 8'h03;
            13'h06CD: rddata <= 8'hCD;
            13'h06CE: rddata <= 8'hA0;
            13'h06CF: rddata <= 8'h0B;
            13'h06D0: rddata <= 8'hC1;
            13'h06D1: rddata <= 8'hE5;
            13'h06D2: rddata <= 8'hE5;
            13'h06D3: rddata <= 8'h2A;
            13'h06D4: rddata <= 8'h4D;
            13'h06D5: rddata <= 8'h38;
            13'h06D6: rddata <= 8'hE3;
            13'h06D7: rddata <= 8'h3E;
            13'h06D8: rddata <= 8'h8C;
            13'h06D9: rddata <= 8'hF5;
            13'h06DA: rddata <= 8'h33;
            13'h06DB: rddata <= 8'hC5;
            13'h06DC: rddata <= 8'hCD;
            13'h06DD: rddata <= 8'h9C;
            13'h06DE: rddata <= 8'h06;
            13'h06DF: rddata <= 8'hCD;
            13'h06E0: rddata <= 8'h1E;
            13'h06E1: rddata <= 8'h07;
            13'h06E2: rddata <= 8'h23;
            13'h06E3: rddata <= 8'hE5;
            13'h06E4: rddata <= 8'h2A;
            13'h06E5: rddata <= 8'h4D;
            13'h06E6: rddata <= 8'h38;
            13'h06E7: rddata <= 8'hE7;
            13'h06E8: rddata <= 8'hE1;
            13'h06E9: rddata <= 8'hDC;
            13'h06EA: rddata <= 8'hA2;
            13'h06EB: rddata <= 8'h04;
            13'h06EC: rddata <= 8'hD4;
            13'h06ED: rddata <= 8'h9F;
            13'h06EE: rddata <= 8'h04;
            13'h06EF: rddata <= 8'h60;
            13'h06F0: rddata <= 8'h69;
            13'h06F1: rddata <= 8'h2B;
            13'h06F2: rddata <= 8'hD8;
            13'h06F3: rddata <= 8'h1E;
            13'h06F4: rddata <= 8'h0E;
            13'h06F5: rddata <= 8'hC3;
            13'h06F6: rddata <= 8'hDB;
            13'h06F7: rddata <= 8'h03;
            13'h06F8: rddata <= 8'hC0;
            13'h06F9: rddata <= 8'h16;
            13'h06FA: rddata <= 8'hFF;
            13'h06FB: rddata <= 8'hCD;
            13'h06FC: rddata <= 8'h9F;
            13'h06FD: rddata <= 8'h03;
            13'h06FE: rddata <= 8'hF9;
            13'h06FF: rddata <= 8'hFE;
            13'h0700: rddata <= 8'h8C;
            13'h0701: rddata <= 8'h1E;
            13'h0702: rddata <= 8'h04;
            13'h0703: rddata <= 8'hC2;
            13'h0704: rddata <= 8'hDB;
            13'h0705: rddata <= 8'h03;
            13'h0706: rddata <= 8'hE1;
            13'h0707: rddata <= 8'h22;
            13'h0708: rddata <= 8'h4D;
            13'h0709: rddata <= 8'h38;
            13'h070A: rddata <= 8'h23;
            13'h070B: rddata <= 8'h7C;
            13'h070C: rddata <= 8'hB5;
            13'h070D: rddata <= 8'h20;
            13'h070E: rddata <= 8'h07;
            13'h070F: rddata <= 8'h3A;
            13'h0710: rddata <= 8'hCC;
            13'h0711: rddata <= 8'h38;
            13'h0712: rddata <= 8'hB7;
            13'h0713: rddata <= 8'hC2;
            13'h0714: rddata <= 8'h01;
            13'h0715: rddata <= 8'h04;
            13'h0716: rddata <= 8'h21;
            13'h0717: rddata <= 8'h2C;
            13'h0718: rddata <= 8'h06;
            13'h0719: rddata <= 8'hE3;
            13'h071A: rddata <= 8'h3E;
            13'h071B: rddata <= 8'hE1;
            13'h071C: rddata <= 8'h01;
            13'h071D: rddata <= 8'h3A;
            13'h071E: rddata <= 8'h0E;
            13'h071F: rddata <= 8'h00;
            13'h0720: rddata <= 8'h06;
            13'h0721: rddata <= 8'h00;
            13'h0722: rddata <= 8'h79;
            13'h0723: rddata <= 8'h48;
            13'h0724: rddata <= 8'h47;
            13'h0725: rddata <= 8'h7E;
            13'h0726: rddata <= 8'hB7;
            13'h0727: rddata <= 8'hC8;
            13'h0728: rddata <= 8'hB8;
            13'h0729: rddata <= 8'hC8;
            13'h072A: rddata <= 8'h23;
            13'h072B: rddata <= 8'hFE;
            13'h072C: rddata <= 8'h22;
            13'h072D: rddata <= 8'h28;
            13'h072E: rddata <= 8'hF3;
            13'h072F: rddata <= 8'h18;
            13'h0730: rddata <= 8'hF4;
            13'h0731: rddata <= 8'hCD;
            13'h0732: rddata <= 8'hD1;
            13'h0733: rddata <= 8'h10;
            13'h0734: rddata <= 8'hCF;
            13'h0735: rddata <= 8'hB0;
            13'h0736: rddata <= 8'hD5;
            13'h0737: rddata <= 8'h3A;
            13'h0738: rddata <= 8'hAB;
            13'h0739: rddata <= 8'h38;
            13'h073A: rddata <= 8'hF5;
            13'h073B: rddata <= 8'hCD;
            13'h073C: rddata <= 8'h85;
            13'h073D: rddata <= 8'h09;
            13'h073E: rddata <= 8'hF1;
            13'h073F: rddata <= 8'hE3;
            13'h0740: rddata <= 8'h22;
            13'h0741: rddata <= 8'hCE;
            13'h0742: rddata <= 8'h38;
            13'h0743: rddata <= 8'h1F;
            13'h0744: rddata <= 8'hCD;
            13'h0745: rddata <= 8'h77;
            13'h0746: rddata <= 8'h09;
            13'h0747: rddata <= 8'hCA;
            13'h0748: rddata <= 8'h79;
            13'h0749: rddata <= 8'h07;
            13'h074A: rddata <= 8'hE5;
            13'h074B: rddata <= 8'h2A;
            13'h074C: rddata <= 8'hE4;
            13'h074D: rddata <= 8'h38;
            13'h074E: rddata <= 8'hE5;
            13'h074F: rddata <= 8'h23;
            13'h0750: rddata <= 8'h23;
            13'h0751: rddata <= 8'h5E;
            13'h0752: rddata <= 8'h23;
            13'h0753: rddata <= 8'h56;
            13'h0754: rddata <= 8'h2A;
            13'h0755: rddata <= 8'h4F;
            13'h0756: rddata <= 8'h38;
            13'h0757: rddata <= 8'hE7;
            13'h0758: rddata <= 8'h30;
            13'h0759: rddata <= 8'h0E;
            13'h075A: rddata <= 8'h2A;
            13'h075B: rddata <= 8'hDA;
            13'h075C: rddata <= 8'h38;
            13'h075D: rddata <= 8'hE7;
            13'h075E: rddata <= 8'hD1;
            13'h075F: rddata <= 8'h30;
            13'h0760: rddata <= 8'h0F;
            13'h0761: rddata <= 8'h21;
            13'h0762: rddata <= 8'hBD;
            13'h0763: rddata <= 8'h38;
            13'h0764: rddata <= 8'hE7;
            13'h0765: rddata <= 8'h30;
            13'h0766: rddata <= 8'h09;
            13'h0767: rddata <= 8'h3E;
            13'h0768: rddata <= 8'hD1;
            13'h0769: rddata <= 8'hCD;
            13'h076A: rddata <= 8'hE4;
            13'h076B: rddata <= 8'h0F;
            13'h076C: rddata <= 8'hEB;
            13'h076D: rddata <= 8'hCD;
            13'h076E: rddata <= 8'h39;
            13'h076F: rddata <= 8'h0E;
            13'h0770: rddata <= 8'hCD;
            13'h0771: rddata <= 8'hE4;
            13'h0772: rddata <= 8'h0F;
            13'h0773: rddata <= 8'hE1;
            13'h0774: rddata <= 8'hCD;
            13'h0775: rddata <= 8'h3D;
            13'h0776: rddata <= 8'h15;
            13'h0777: rddata <= 8'hE1;
            13'h0778: rddata <= 8'hC9;
            13'h0779: rddata <= 8'hE5;
            13'h077A: rddata <= 8'hCD;
            13'h077B: rddata <= 8'h3A;
            13'h077C: rddata <= 8'h15;
            13'h077D: rddata <= 8'hD1;
            13'h077E: rddata <= 8'hE1;
            13'h077F: rddata <= 8'hC9;
            13'h0780: rddata <= 8'hF7;
            13'h0781: rddata <= 8'h19;
            13'h0782: rddata <= 8'hCD;
            13'h0783: rddata <= 8'h54;
            13'h0784: rddata <= 8'h0B;
            13'h0785: rddata <= 8'h7E;
            13'h0786: rddata <= 8'h47;
            13'h0787: rddata <= 8'hFE;
            13'h0788: rddata <= 8'h8C;
            13'h0789: rddata <= 8'h28;
            13'h078A: rddata <= 8'h03;
            13'h078B: rddata <= 8'hCF;
            13'h078C: rddata <= 8'h88;
            13'h078D: rddata <= 8'h2B;
            13'h078E: rddata <= 8'h4B;
            13'h078F: rddata <= 8'h0D;
            13'h0790: rddata <= 8'h78;
            13'h0791: rddata <= 8'hCA;
            13'h0792: rddata <= 8'h51;
            13'h0793: rddata <= 8'h06;
            13'h0794: rddata <= 8'hCD;
            13'h0795: rddata <= 8'h9D;
            13'h0796: rddata <= 8'h06;
            13'h0797: rddata <= 8'hFE;
            13'h0798: rddata <= 8'h2C;
            13'h0799: rddata <= 8'hC0;
            13'h079A: rddata <= 8'h18;
            13'h079B: rddata <= 8'hF3;
            13'h079C: rddata <= 8'hCD;
            13'h079D: rddata <= 8'h85;
            13'h079E: rddata <= 8'h09;
            13'h079F: rddata <= 8'h7E;
            13'h07A0: rddata <= 8'hFE;
            13'h07A1: rddata <= 8'h88;
            13'h07A2: rddata <= 8'h28;
            13'h07A3: rddata <= 8'h03;
            13'h07A4: rddata <= 8'hCF;
            13'h07A5: rddata <= 8'hA5;
            13'h07A6: rddata <= 8'h2B;
            13'h07A7: rddata <= 8'hCD;
            13'h07A8: rddata <= 8'h75;
            13'h07A9: rddata <= 8'h09;
            13'h07AA: rddata <= 8'hEF;
            13'h07AB: rddata <= 8'hCA;
            13'h07AC: rddata <= 8'h1E;
            13'h07AD: rddata <= 8'h07;
            13'h07AE: rddata <= 8'hD7;
            13'h07AF: rddata <= 8'hDA;
            13'h07B0: rddata <= 8'hDC;
            13'h07B1: rddata <= 8'h06;
            13'h07B2: rddata <= 8'hC3;
            13'h07B3: rddata <= 8'h50;
            13'h07B4: rddata <= 8'h06;
            13'h07B5: rddata <= 8'h3E;
            13'h07B6: rddata <= 8'h01;
            13'h07B7: rddata <= 8'h32;
            13'h07B8: rddata <= 8'h47;
            13'h07B9: rddata <= 8'h38;
            13'h07BA: rddata <= 8'h2B;
            13'h07BB: rddata <= 8'hD7;
            13'h07BC: rddata <= 8'hF7;
            13'h07BD: rddata <= 8'h06;
            13'h07BE: rddata <= 8'hCC;
            13'h07BF: rddata <= 8'hEA;
            13'h07C0: rddata <= 8'h19;
            13'h07C1: rddata <= 8'hCA;
            13'h07C2: rddata <= 8'h66;
            13'h07C3: rddata <= 8'h08;
            13'h07C4: rddata <= 8'hFE;
            13'h07C5: rddata <= 8'hA0;
            13'h07C6: rddata <= 8'hCA;
            13'h07C7: rddata <= 8'h3A;
            13'h07C8: rddata <= 8'h08;
            13'h07C9: rddata <= 8'hFE;
            13'h07CA: rddata <= 8'hA3;
            13'h07CB: rddata <= 8'hCA;
            13'h07CC: rddata <= 8'h3A;
            13'h07CD: rddata <= 8'h08;
            13'h07CE: rddata <= 8'hE5;
            13'h07CF: rddata <= 8'hFE;
            13'h07D0: rddata <= 8'h2C;
            13'h07D1: rddata <= 8'h28;
            13'h07D2: rddata <= 8'h44;
            13'h07D3: rddata <= 8'hFE;
            13'h07D4: rddata <= 8'h3B;
            13'h07D5: rddata <= 8'hCA;
            13'h07D6: rddata <= 8'h61;
            13'h07D7: rddata <= 8'h08;
            13'h07D8: rddata <= 8'hC1;
            13'h07D9: rddata <= 8'hCD;
            13'h07DA: rddata <= 8'h85;
            13'h07DB: rddata <= 8'h09;
            13'h07DC: rddata <= 8'hE5;
            13'h07DD: rddata <= 8'h3A;
            13'h07DE: rddata <= 8'hAB;
            13'h07DF: rddata <= 8'h38;
            13'h07E0: rddata <= 8'hB7;
            13'h07E1: rddata <= 8'hC2;
            13'h07E2: rddata <= 8'h11;
            13'h07E3: rddata <= 8'h08;
            13'h07E4: rddata <= 8'hCD;
            13'h07E5: rddata <= 8'h80;
            13'h07E6: rddata <= 8'h16;
            13'h07E7: rddata <= 8'hCD;
            13'h07E8: rddata <= 8'h5F;
            13'h07E9: rddata <= 8'h0E;
            13'h07EA: rddata <= 8'h36;
            13'h07EB: rddata <= 8'h20;
            13'h07EC: rddata <= 8'h2A;
            13'h07ED: rddata <= 8'hE4;
            13'h07EE: rddata <= 8'h38;
            13'h07EF: rddata <= 8'h3A;
            13'h07F0: rddata <= 8'h47;
            13'h07F1: rddata <= 8'h38;
            13'h07F2: rddata <= 8'hB7;
            13'h07F3: rddata <= 8'h28;
            13'h07F4: rddata <= 8'h08;
            13'h07F5: rddata <= 8'h3A;
            13'h07F6: rddata <= 8'h46;
            13'h07F7: rddata <= 8'h38;
            13'h07F8: rddata <= 8'h86;
            13'h07F9: rddata <= 8'hFE;
            13'h07FA: rddata <= 8'h84;
            13'h07FB: rddata <= 8'h18;
            13'h07FC: rddata <= 8'h0D;
            13'h07FD: rddata <= 8'h3A;
            13'h07FE: rddata <= 8'h48;
            13'h07FF: rddata <= 8'h38;
            13'h0800: rddata <= 8'h47;
            13'h0801: rddata <= 8'h3C;
            13'h0802: rddata <= 8'h28;
            13'h0803: rddata <= 8'h09;
            13'h0804: rddata <= 8'h3A;
            13'h0805: rddata <= 8'h00;
            13'h0806: rddata <= 8'h38;
            13'h0807: rddata <= 8'h86;
            13'h0808: rddata <= 8'h3D;
            13'h0809: rddata <= 8'hB8;
            13'h080A: rddata <= 8'hD4;
            13'h080B: rddata <= 8'hEA;
            13'h080C: rddata <= 8'h19;
            13'h080D: rddata <= 8'hCD;
            13'h080E: rddata <= 8'hA0;
            13'h080F: rddata <= 8'h0E;
            13'h0810: rddata <= 8'hAF;
            13'h0811: rddata <= 8'hC4;
            13'h0812: rddata <= 8'hA0;
            13'h0813: rddata <= 8'h0E;
            13'h0814: rddata <= 8'hE1;
            13'h0815: rddata <= 8'h18;
            13'h0816: rddata <= 8'hA3;
            13'h0817: rddata <= 8'h3A;
            13'h0818: rddata <= 8'h47;
            13'h0819: rddata <= 8'h38;
            13'h081A: rddata <= 8'hB7;
            13'h081B: rddata <= 8'h28;
            13'h081C: rddata <= 8'h08;
            13'h081D: rddata <= 8'h3A;
            13'h081E: rddata <= 8'h46;
            13'h081F: rddata <= 8'h38;
            13'h0820: rddata <= 8'hFE;
            13'h0821: rddata <= 8'h70;
            13'h0822: rddata <= 8'hC3;
            13'h0823: rddata <= 8'h2D;
            13'h0824: rddata <= 8'h08;
            13'h0825: rddata <= 8'h3A;
            13'h0826: rddata <= 8'h49;
            13'h0827: rddata <= 8'h38;
            13'h0828: rddata <= 8'h47;
            13'h0829: rddata <= 8'h3A;
            13'h082A: rddata <= 8'h00;
            13'h082B: rddata <= 8'h38;
            13'h082C: rddata <= 8'hB8;
            13'h082D: rddata <= 8'hD4;
            13'h082E: rddata <= 8'hEA;
            13'h082F: rddata <= 8'h19;
            13'h0830: rddata <= 8'hD2;
            13'h0831: rddata <= 8'h61;
            13'h0832: rddata <= 8'h08;
            13'h0833: rddata <= 8'hD6;
            13'h0834: rddata <= 8'h0E;
            13'h0835: rddata <= 8'h30;
            13'h0836: rddata <= 8'hFC;
            13'h0837: rddata <= 8'h2F;
            13'h0838: rddata <= 8'h18;
            13'h0839: rddata <= 8'h20;
            13'h083A: rddata <= 8'hF5;
            13'h083B: rddata <= 8'hCD;
            13'h083C: rddata <= 8'h53;
            13'h083D: rddata <= 8'h0B;
            13'h083E: rddata <= 8'hCF;
            13'h083F: rddata <= 8'h29;
            13'h0840: rddata <= 8'h2B;
            13'h0841: rddata <= 8'hF1;
            13'h0842: rddata <= 8'hD6;
            13'h0843: rddata <= 8'hA3;
            13'h0844: rddata <= 8'hE5;
            13'h0845: rddata <= 8'h28;
            13'h0846: rddata <= 8'h0F;
            13'h0847: rddata <= 8'h3A;
            13'h0848: rddata <= 8'h47;
            13'h0849: rddata <= 8'h38;
            13'h084A: rddata <= 8'hB7;
            13'h084B: rddata <= 8'hCA;
            13'h084C: rddata <= 8'h53;
            13'h084D: rddata <= 8'h08;
            13'h084E: rddata <= 8'h3A;
            13'h084F: rddata <= 8'h46;
            13'h0850: rddata <= 8'h38;
            13'h0851: rddata <= 8'h18;
            13'h0852: rddata <= 8'h03;
            13'h0853: rddata <= 8'h3A;
            13'h0854: rddata <= 8'h00;
            13'h0855: rddata <= 8'h38;
            13'h0856: rddata <= 8'h2F;
            13'h0857: rddata <= 8'h83;
            13'h0858: rddata <= 8'h30;
            13'h0859: rddata <= 8'h07;
            13'h085A: rddata <= 8'h3C;
            13'h085B: rddata <= 8'h47;
            13'h085C: rddata <= 8'h3E;
            13'h085D: rddata <= 8'h20;
            13'h085E: rddata <= 8'hDF;
            13'h085F: rddata <= 8'h10;
            13'h0860: rddata <= 8'hFD;
            13'h0861: rddata <= 8'hE1;
            13'h0862: rddata <= 8'hD7;
            13'h0863: rddata <= 8'hC3;
            13'h0864: rddata <= 8'hC1;
            13'h0865: rddata <= 8'h07;
            13'h0866: rddata <= 8'hF7;
            13'h0867: rddata <= 8'h07;
            13'h0868: rddata <= 8'hAF;
            13'h0869: rddata <= 8'h32;
            13'h086A: rddata <= 8'h47;
            13'h086B: rddata <= 8'h38;
            13'h086C: rddata <= 8'hC9;
            13'h086D: rddata <= 8'h3F;
            13'h086E: rddata <= 8'h52;
            13'h086F: rddata <= 8'h65;
            13'h0870: rddata <= 8'h64;
            13'h0871: rddata <= 8'h6F;
            13'h0872: rddata <= 8'h20;
            13'h0873: rddata <= 8'h66;
            13'h0874: rddata <= 8'h72;
            13'h0875: rddata <= 8'h6F;
            13'h0876: rddata <= 8'h6D;
            13'h0877: rddata <= 8'h20;
            13'h0878: rddata <= 8'h73;
            13'h0879: rddata <= 8'h74;
            13'h087A: rddata <= 8'h61;
            13'h087B: rddata <= 8'h72;
            13'h087C: rddata <= 8'h74;
            13'h087D: rddata <= 8'h0D;
            13'h087E: rddata <= 8'h0A;
            13'h087F: rddata <= 8'h00;
            13'h0880: rddata <= 8'hF7;
            13'h0881: rddata <= 8'h08;
            13'h0882: rddata <= 8'h3A;
            13'h0883: rddata <= 8'hCD;
            13'h0884: rddata <= 8'h38;
            13'h0885: rddata <= 8'hB7;
            13'h0886: rddata <= 8'hC2;
            13'h0887: rddata <= 8'hBE;
            13'h0888: rddata <= 8'h03;
            13'h0889: rddata <= 8'hC1;
            13'h088A: rddata <= 8'h21;
            13'h088B: rddata <= 8'h6D;
            13'h088C: rddata <= 8'h08;
            13'h088D: rddata <= 8'hCD;
            13'h088E: rddata <= 8'h9D;
            13'h088F: rddata <= 8'h0E;
            13'h0890: rddata <= 8'hC3;
            13'h0891: rddata <= 8'h01;
            13'h0892: rddata <= 8'h0C;
            13'h0893: rddata <= 8'hF7;
            13'h0894: rddata <= 8'h1A;
            13'h0895: rddata <= 8'hCD;
            13'h0896: rddata <= 8'h45;
            13'h0897: rddata <= 8'h0B;
            13'h0898: rddata <= 8'h7E;
            13'h0899: rddata <= 8'hFE;
            13'h089A: rddata <= 8'h22;
            13'h089B: rddata <= 8'h3E;
            13'h089C: rddata <= 8'h00;
            13'h089D: rddata <= 8'hC2;
            13'h089E: rddata <= 8'hAA;
            13'h089F: rddata <= 8'h08;
            13'h08A0: rddata <= 8'hCD;
            13'h08A1: rddata <= 8'h60;
            13'h08A2: rddata <= 8'h0E;
            13'h08A3: rddata <= 8'hCF;
            13'h08A4: rddata <= 8'h3B;
            13'h08A5: rddata <= 8'hE5;
            13'h08A6: rddata <= 8'hCD;
            13'h08A7: rddata <= 8'hA0;
            13'h08A8: rddata <= 8'h0E;
            13'h08A9: rddata <= 8'h3E;
            13'h08AA: rddata <= 8'hE5;
            13'h08AB: rddata <= 8'hCD;
            13'h08AC: rddata <= 8'h5B;
            13'h08AD: rddata <= 8'h0D;
            13'h08AE: rddata <= 8'hC1;
            13'h08AF: rddata <= 8'hDA;
            13'h08B0: rddata <= 8'h26;
            13'h08B1: rddata <= 8'h0C;
            13'h08B2: rddata <= 8'h23;
            13'h08B3: rddata <= 8'h7E;
            13'h08B4: rddata <= 8'hB7;
            13'h08B5: rddata <= 8'h2B;
            13'h08B6: rddata <= 8'hC5;
            13'h08B7: rddata <= 8'hCA;
            13'h08B8: rddata <= 8'h1B;
            13'h08B9: rddata <= 8'h07;
            13'h08BA: rddata <= 8'h36;
            13'h08BB: rddata <= 8'h2C;
            13'h08BC: rddata <= 8'h18;
            13'h08BD: rddata <= 8'h05;
            13'h08BE: rddata <= 8'hE5;
            13'h08BF: rddata <= 8'h2A;
            13'h08C0: rddata <= 8'hDC;
            13'h08C1: rddata <= 8'h38;
            13'h08C2: rddata <= 8'hF6;
            13'h08C3: rddata <= 8'hAF;
            13'h08C4: rddata <= 8'h32;
            13'h08C5: rddata <= 8'hCD;
            13'h08C6: rddata <= 8'h38;
            13'h08C7: rddata <= 8'hE3;
            13'h08C8: rddata <= 8'h01;
            13'h08C9: rddata <= 8'hCF;
            13'h08CA: rddata <= 8'h2C;
            13'h08CB: rddata <= 8'hCD;
            13'h08CC: rddata <= 8'hD1;
            13'h08CD: rddata <= 8'h10;
            13'h08CE: rddata <= 8'hE3;
            13'h08CF: rddata <= 8'hD5;
            13'h08D0: rddata <= 8'h7E;
            13'h08D1: rddata <= 8'hFE;
            13'h08D2: rddata <= 8'h2C;
            13'h08D3: rddata <= 8'h28;
            13'h08D4: rddata <= 8'h1B;
            13'h08D5: rddata <= 8'h3A;
            13'h08D6: rddata <= 8'hCD;
            13'h08D7: rddata <= 8'h38;
            13'h08D8: rddata <= 8'hB7;
            13'h08D9: rddata <= 8'hC2;
            13'h08DA: rddata <= 8'h53;
            13'h08DB: rddata <= 8'h09;
            13'h08DC: rddata <= 8'h3E;
            13'h08DD: rddata <= 8'h3F;
            13'h08DE: rddata <= 8'hDF;
            13'h08DF: rddata <= 8'hCD;
            13'h08E0: rddata <= 8'h5B;
            13'h08E1: rddata <= 8'h0D;
            13'h08E2: rddata <= 8'hD1;
            13'h08E3: rddata <= 8'hC1;
            13'h08E4: rddata <= 8'hDA;
            13'h08E5: rddata <= 8'h26;
            13'h08E6: rddata <= 8'h0C;
            13'h08E7: rddata <= 8'h23;
            13'h08E8: rddata <= 8'h7E;
            13'h08E9: rddata <= 8'h2B;
            13'h08EA: rddata <= 8'hB7;
            13'h08EB: rddata <= 8'hC5;
            13'h08EC: rddata <= 8'hCA;
            13'h08ED: rddata <= 8'h1B;
            13'h08EE: rddata <= 8'h07;
            13'h08EF: rddata <= 8'hD5;
            13'h08F0: rddata <= 8'hF7;
            13'h08F1: rddata <= 8'h1C;
            13'h08F2: rddata <= 8'h3A;
            13'h08F3: rddata <= 8'hAB;
            13'h08F4: rddata <= 8'h38;
            13'h08F5: rddata <= 8'hB7;
            13'h08F6: rddata <= 8'h28;
            13'h08F7: rddata <= 8'h1F;
            13'h08F8: rddata <= 8'hD7;
            13'h08F9: rddata <= 8'h57;
            13'h08FA: rddata <= 8'h47;
            13'h08FB: rddata <= 8'hFE;
            13'h08FC: rddata <= 8'h22;
            13'h08FD: rddata <= 8'h28;
            13'h08FE: rddata <= 8'h0C;
            13'h08FF: rddata <= 8'h3A;
            13'h0900: rddata <= 8'hCD;
            13'h0901: rddata <= 8'h38;
            13'h0902: rddata <= 8'hB7;
            13'h0903: rddata <= 8'h57;
            13'h0904: rddata <= 8'h28;
            13'h0905: rddata <= 8'h02;
            13'h0906: rddata <= 8'h16;
            13'h0907: rddata <= 8'h3A;
            13'h0908: rddata <= 8'h06;
            13'h0909: rddata <= 8'h2C;
            13'h090A: rddata <= 8'h2B;
            13'h090B: rddata <= 8'hCD;
            13'h090C: rddata <= 8'h63;
            13'h090D: rddata <= 8'h0E;
            13'h090E: rddata <= 8'hEB;
            13'h090F: rddata <= 8'h21;
            13'h0910: rddata <= 8'h20;
            13'h0911: rddata <= 8'h09;
            13'h0912: rddata <= 8'hE3;
            13'h0913: rddata <= 8'hD5;
            13'h0914: rddata <= 8'hC3;
            13'h0915: rddata <= 8'h4A;
            13'h0916: rddata <= 8'h07;
            13'h0917: rddata <= 8'hD7;
            13'h0918: rddata <= 8'hCD;
            13'h0919: rddata <= 8'hE5;
            13'h091A: rddata <= 8'h15;
            13'h091B: rddata <= 8'hE3;
            13'h091C: rddata <= 8'hCD;
            13'h091D: rddata <= 8'h3A;
            13'h091E: rddata <= 8'h15;
            13'h091F: rddata <= 8'hE1;
            13'h0920: rddata <= 8'h2B;
            13'h0921: rddata <= 8'hD7;
            13'h0922: rddata <= 8'h28;
            13'h0923: rddata <= 8'h05;
            13'h0924: rddata <= 8'hFE;
            13'h0925: rddata <= 8'h2C;
            13'h0926: rddata <= 8'hC2;
            13'h0927: rddata <= 8'h80;
            13'h0928: rddata <= 8'h08;
            13'h0929: rddata <= 8'hE3;
            13'h092A: rddata <= 8'h2B;
            13'h092B: rddata <= 8'hD7;
            13'h092C: rddata <= 8'hC2;
            13'h092D: rddata <= 8'hC9;
            13'h092E: rddata <= 8'h08;
            13'h092F: rddata <= 8'hD1;
            13'h0930: rddata <= 8'h3A;
            13'h0931: rddata <= 8'hCD;
            13'h0932: rddata <= 8'h38;
            13'h0933: rddata <= 8'hB7;
            13'h0934: rddata <= 8'hEB;
            13'h0935: rddata <= 8'hC2;
            13'h0936: rddata <= 8'h1A;
            13'h0937: rddata <= 8'h0C;
            13'h0938: rddata <= 8'hD5;
            13'h0939: rddata <= 8'hB6;
            13'h093A: rddata <= 8'h21;
            13'h093B: rddata <= 8'h42;
            13'h093C: rddata <= 8'h09;
            13'h093D: rddata <= 8'hC4;
            13'h093E: rddata <= 8'h9D;
            13'h093F: rddata <= 8'h0E;
            13'h0940: rddata <= 8'hE1;
            13'h0941: rddata <= 8'hC9;
            13'h0942: rddata <= 8'h3F;
            13'h0943: rddata <= 8'h45;
            13'h0944: rddata <= 8'h78;
            13'h0945: rddata <= 8'h74;
            13'h0946: rddata <= 8'h72;
            13'h0947: rddata <= 8'h61;
            13'h0948: rddata <= 8'h20;
            13'h0949: rddata <= 8'h69;
            13'h094A: rddata <= 8'h67;
            13'h094B: rddata <= 8'h6E;
            13'h094C: rddata <= 8'h6F;
            13'h094D: rddata <= 8'h72;
            13'h094E: rddata <= 8'h65;
            13'h094F: rddata <= 8'h64;
            13'h0950: rddata <= 8'h0D;
            13'h0951: rddata <= 8'h0A;
            13'h0952: rddata <= 8'h00;
            13'h0953: rddata <= 8'hCD;
            13'h0954: rddata <= 8'h1C;
            13'h0955: rddata <= 8'h07;
            13'h0956: rddata <= 8'hB7;
            13'h0957: rddata <= 8'h20;
            13'h0958: rddata <= 8'h11;
            13'h0959: rddata <= 8'h23;
            13'h095A: rddata <= 8'h7E;
            13'h095B: rddata <= 8'h23;
            13'h095C: rddata <= 8'hB6;
            13'h095D: rddata <= 8'h1E;
            13'h095E: rddata <= 8'h06;
            13'h095F: rddata <= 8'hCA;
            13'h0960: rddata <= 8'hDB;
            13'h0961: rddata <= 8'h03;
            13'h0962: rddata <= 8'h23;
            13'h0963: rddata <= 8'h5E;
            13'h0964: rddata <= 8'h23;
            13'h0965: rddata <= 8'h56;
            13'h0966: rddata <= 8'hED;
            13'h0967: rddata <= 8'h53;
            13'h0968: rddata <= 8'hC9;
            13'h0969: rddata <= 8'h38;
            13'h096A: rddata <= 8'hD7;
            13'h096B: rddata <= 8'hFE;
            13'h096C: rddata <= 8'h83;
            13'h096D: rddata <= 8'h20;
            13'h096E: rddata <= 8'hE4;
            13'h096F: rddata <= 8'hC3;
            13'h0970: rddata <= 8'hF0;
            13'h0971: rddata <= 8'h08;
            13'h0972: rddata <= 8'hCD;
            13'h0973: rddata <= 8'h85;
            13'h0974: rddata <= 8'h09;
            13'h0975: rddata <= 8'hF6;
            13'h0976: rddata <= 8'h37;
            13'h0977: rddata <= 8'h3A;
            13'h0978: rddata <= 8'hAB;
            13'h0979: rddata <= 8'h38;
            13'h097A: rddata <= 8'h8F;
            13'h097B: rddata <= 8'hB7;
            13'h097C: rddata <= 8'hE8;
            13'h097D: rddata <= 8'hC3;
            13'h097E: rddata <= 8'hD9;
            13'h097F: rddata <= 8'h03;
            13'h0980: rddata <= 8'hCF;
            13'h0981: rddata <= 8'hB0;
            13'h0982: rddata <= 8'h01;
            13'h0983: rddata <= 8'hCF;
            13'h0984: rddata <= 8'h28;
            13'h0985: rddata <= 8'h2B;
            13'h0986: rddata <= 8'h16;
            13'h0987: rddata <= 8'h00;
            13'h0988: rddata <= 8'hD5;
            13'h0989: rddata <= 8'h0E;
            13'h098A: rddata <= 8'h01;
            13'h098B: rddata <= 8'hCD;
            13'h098C: rddata <= 8'hA0;
            13'h098D: rddata <= 8'h0B;
            13'h098E: rddata <= 8'hCD;
            13'h098F: rddata <= 8'hFD;
            13'h0990: rddata <= 8'h09;
            13'h0991: rddata <= 8'h22;
            13'h0992: rddata <= 8'hD0;
            13'h0993: rddata <= 8'h38;
            13'h0994: rddata <= 8'h2A;
            13'h0995: rddata <= 8'hD0;
            13'h0996: rddata <= 8'h38;
            13'h0997: rddata <= 8'hC1;
            13'h0998: rddata <= 8'h78;
            13'h0999: rddata <= 8'hFE;
            13'h099A: rddata <= 8'h78;
            13'h099B: rddata <= 8'hD4;
            13'h099C: rddata <= 8'h75;
            13'h099D: rddata <= 8'h09;
            13'h099E: rddata <= 8'h7E;
            13'h099F: rddata <= 8'h22;
            13'h09A0: rddata <= 8'hC3;
            13'h09A1: rddata <= 8'h38;
            13'h09A2: rddata <= 8'hFE;
            13'h09A3: rddata <= 8'hA8;
            13'h09A4: rddata <= 8'hD8;
            13'h09A5: rddata <= 8'hFE;
            13'h09A6: rddata <= 8'hB2;
            13'h09A7: rddata <= 8'hD0;
            13'h09A8: rddata <= 8'hFE;
            13'h09A9: rddata <= 8'hAF;
            13'h09AA: rddata <= 8'hD2;
            13'h09AB: rddata <= 8'hE2;
            13'h09AC: rddata <= 8'h09;
            13'h09AD: rddata <= 8'hD6;
            13'h09AE: rddata <= 8'hA8;
            13'h09AF: rddata <= 8'h5F;
            13'h09B0: rddata <= 8'h20;
            13'h09B1: rddata <= 8'h08;
            13'h09B2: rddata <= 8'h3A;
            13'h09B3: rddata <= 8'hAB;
            13'h09B4: rddata <= 8'h38;
            13'h09B5: rddata <= 8'h3D;
            13'h09B6: rddata <= 8'h7B;
            13'h09B7: rddata <= 8'hCA;
            13'h09B8: rddata <= 8'h7C;
            13'h09B9: rddata <= 8'h0F;
            13'h09BA: rddata <= 8'h07;
            13'h09BB: rddata <= 8'h83;
            13'h09BC: rddata <= 8'h5F;
            13'h09BD: rddata <= 8'h21;
            13'h09BE: rddata <= 8'h4C;
            13'h09BF: rddata <= 8'h03;
            13'h09C0: rddata <= 8'h16;
            13'h09C1: rddata <= 8'h00;
            13'h09C2: rddata <= 8'h19;
            13'h09C3: rddata <= 8'h78;
            13'h09C4: rddata <= 8'h56;
            13'h09C5: rddata <= 8'hBA;
            13'h09C6: rddata <= 8'hD0;
            13'h09C7: rddata <= 8'h23;
            13'h09C8: rddata <= 8'hCD;
            13'h09C9: rddata <= 8'h75;
            13'h09CA: rddata <= 8'h09;
            13'h09CB: rddata <= 8'hC5;
            13'h09CC: rddata <= 8'h01;
            13'h09CD: rddata <= 8'h94;
            13'h09CE: rddata <= 8'h09;
            13'h09CF: rddata <= 8'hC5;
            13'h09D0: rddata <= 8'h43;
            13'h09D1: rddata <= 8'h4A;
            13'h09D2: rddata <= 8'hCD;
            13'h09D3: rddata <= 8'h13;
            13'h09D4: rddata <= 8'h15;
            13'h09D5: rddata <= 8'h58;
            13'h09D6: rddata <= 8'h51;
            13'h09D7: rddata <= 8'h4E;
            13'h09D8: rddata <= 8'h23;
            13'h09D9: rddata <= 8'h46;
            13'h09DA: rddata <= 8'h23;
            13'h09DB: rddata <= 8'hC5;
            13'h09DC: rddata <= 8'h2A;
            13'h09DD: rddata <= 8'hC3;
            13'h09DE: rddata <= 8'h38;
            13'h09DF: rddata <= 8'hC3;
            13'h09E0: rddata <= 8'h88;
            13'h09E1: rddata <= 8'h09;
            13'h09E2: rddata <= 8'h16;
            13'h09E3: rddata <= 8'h00;
            13'h09E4: rddata <= 8'hD6;
            13'h09E5: rddata <= 8'hAF;
            13'h09E6: rddata <= 8'hDA;
            13'h09E7: rddata <= 8'hD0;
            13'h09E8: rddata <= 8'h0A;
            13'h09E9: rddata <= 8'hFE;
            13'h09EA: rddata <= 8'h03;
            13'h09EB: rddata <= 8'hD2;
            13'h09EC: rddata <= 8'hD0;
            13'h09ED: rddata <= 8'h0A;
            13'h09EE: rddata <= 8'hFE;
            13'h09EF: rddata <= 8'h01;
            13'h09F0: rddata <= 8'h17;
            13'h09F1: rddata <= 8'hAA;
            13'h09F2: rddata <= 8'hBA;
            13'h09F3: rddata <= 8'h57;
            13'h09F4: rddata <= 8'hDA;
            13'h09F5: rddata <= 8'hC4;
            13'h09F6: rddata <= 8'h03;
            13'h09F7: rddata <= 8'h22;
            13'h09F8: rddata <= 8'hC3;
            13'h09F9: rddata <= 8'h38;
            13'h09FA: rddata <= 8'hD7;
            13'h09FB: rddata <= 8'h18;
            13'h09FC: rddata <= 8'hE7;
            13'h09FD: rddata <= 8'hF7;
            13'h09FE: rddata <= 8'h09;
            13'h09FF: rddata <= 8'hAF;
            13'h0A00: rddata <= 8'h32;
            13'h0A01: rddata <= 8'hAB;
            13'h0A02: rddata <= 8'h38;
            13'h0A03: rddata <= 8'hD7;
            13'h0A04: rddata <= 8'hCA;
            13'h0A05: rddata <= 8'hD6;
            13'h0A06: rddata <= 8'h03;
            13'h0A07: rddata <= 8'hDA;
            13'h0A08: rddata <= 8'hE5;
            13'h0A09: rddata <= 8'h15;
            13'h0A0A: rddata <= 8'hCD;
            13'h0A0B: rddata <= 8'hC6;
            13'h0A0C: rddata <= 8'h0C;
            13'h0A0D: rddata <= 8'hD2;
            13'h0A0E: rddata <= 8'h4E;
            13'h0A0F: rddata <= 8'h0A;
            13'h0A10: rddata <= 8'hFE;
            13'h0A11: rddata <= 8'hA8;
            13'h0A12: rddata <= 8'h28;
            13'h0A13: rddata <= 8'hE9;
            13'h0A14: rddata <= 8'hFE;
            13'h0A15: rddata <= 8'h2E;
            13'h0A16: rddata <= 8'hCA;
            13'h0A17: rddata <= 8'hE5;
            13'h0A18: rddata <= 8'h15;
            13'h0A19: rddata <= 8'hFE;
            13'h0A1A: rddata <= 8'hA9;
            13'h0A1B: rddata <= 8'hCA;
            13'h0A1C: rddata <= 8'h3D;
            13'h0A1D: rddata <= 8'h0A;
            13'h0A1E: rddata <= 8'hFE;
            13'h0A1F: rddata <= 8'h22;
            13'h0A20: rddata <= 8'hCA;
            13'h0A21: rddata <= 8'h60;
            13'h0A22: rddata <= 8'h0E;
            13'h0A23: rddata <= 8'hFE;
            13'h0A24: rddata <= 8'hA6;
            13'h0A25: rddata <= 8'hCA;
            13'h0A26: rddata <= 8'h05;
            13'h0A27: rddata <= 8'h0B;
            13'h0A28: rddata <= 8'hFE;
            13'h0A29: rddata <= 8'hA4;
            13'h0A2A: rddata <= 8'hCA;
            13'h0A2B: rddata <= 8'hFB;
            13'h0A2C: rddata <= 8'h19;
            13'h0A2D: rddata <= 8'hFE;
            13'h0A2E: rddata <= 8'hA2;
            13'h0A2F: rddata <= 8'hCA;
            13'h0A30: rddata <= 8'h40;
            13'h0A31: rddata <= 8'h0B;
            13'h0A32: rddata <= 8'hD6;
            13'h0A33: rddata <= 8'hB2;
            13'h0A34: rddata <= 8'hD2;
            13'h0A35: rddata <= 8'h5F;
            13'h0A36: rddata <= 8'h0A;
            13'h0A37: rddata <= 8'hCD;
            13'h0A38: rddata <= 8'h83;
            13'h0A39: rddata <= 8'h09;
            13'h0A3A: rddata <= 8'hCF;
            13'h0A3B: rddata <= 8'h29;
            13'h0A3C: rddata <= 8'hC9;
            13'h0A3D: rddata <= 8'h16;
            13'h0A3E: rddata <= 8'h7D;
            13'h0A3F: rddata <= 8'hCD;
            13'h0A40: rddata <= 8'h88;
            13'h0A41: rddata <= 8'h09;
            13'h0A42: rddata <= 8'h2A;
            13'h0A43: rddata <= 8'hD0;
            13'h0A44: rddata <= 8'h38;
            13'h0A45: rddata <= 8'hE5;
            13'h0A46: rddata <= 8'hCD;
            13'h0A47: rddata <= 8'h0B;
            13'h0A48: rddata <= 8'h15;
            13'h0A49: rddata <= 8'hCD;
            13'h0A4A: rddata <= 8'h75;
            13'h0A4B: rddata <= 8'h09;
            13'h0A4C: rddata <= 8'hE1;
            13'h0A4D: rddata <= 8'hC9;
            13'h0A4E: rddata <= 8'hCD;
            13'h0A4F: rddata <= 8'hD1;
            13'h0A50: rddata <= 8'h10;
            13'h0A51: rddata <= 8'hE5;
            13'h0A52: rddata <= 8'hEB;
            13'h0A53: rddata <= 8'h22;
            13'h0A54: rddata <= 8'hE4;
            13'h0A55: rddata <= 8'h38;
            13'h0A56: rddata <= 8'h3A;
            13'h0A57: rddata <= 8'hAB;
            13'h0A58: rddata <= 8'h38;
            13'h0A59: rddata <= 8'hB7;
            13'h0A5A: rddata <= 8'hCC;
            13'h0A5B: rddata <= 8'h20;
            13'h0A5C: rddata <= 8'h15;
            13'h0A5D: rddata <= 8'hE1;
            13'h0A5E: rddata <= 8'hC9;
            13'h0A5F: rddata <= 8'hF7;
            13'h0A60: rddata <= 8'h1B;
            13'h0A61: rddata <= 8'hFE;
            13'h0A62: rddata <= 8'h18;
            13'h0A63: rddata <= 8'hCA;
            13'h0A64: rddata <= 8'h68;
            13'h0A65: rddata <= 8'h1A;
            13'h0A66: rddata <= 8'h06;
            13'h0A67: rddata <= 8'h00;
            13'h0A68: rddata <= 8'h07;
            13'h0A69: rddata <= 8'h4F;
            13'h0A6A: rddata <= 8'hC5;
            13'h0A6B: rddata <= 8'hD7;
            13'h0A6C: rddata <= 8'h79;
            13'h0A6D: rddata <= 8'hFE;
            13'h0A6E: rddata <= 8'h29;
            13'h0A6F: rddata <= 8'h38;
            13'h0A70: rddata <= 8'h16;
            13'h0A71: rddata <= 8'hCD;
            13'h0A72: rddata <= 8'h83;
            13'h0A73: rddata <= 8'h09;
            13'h0A74: rddata <= 8'hCF;
            13'h0A75: rddata <= 8'h2C;
            13'h0A76: rddata <= 8'hCD;
            13'h0A77: rddata <= 8'h76;
            13'h0A78: rddata <= 8'h09;
            13'h0A79: rddata <= 8'hEB;
            13'h0A7A: rddata <= 8'h2A;
            13'h0A7B: rddata <= 8'hE4;
            13'h0A7C: rddata <= 8'h38;
            13'h0A7D: rddata <= 8'hE3;
            13'h0A7E: rddata <= 8'hE5;
            13'h0A7F: rddata <= 8'hEB;
            13'h0A80: rddata <= 8'hCD;
            13'h0A81: rddata <= 8'h54;
            13'h0A82: rddata <= 8'h0B;
            13'h0A83: rddata <= 8'hEB;
            13'h0A84: rddata <= 8'hE3;
            13'h0A85: rddata <= 8'h18;
            13'h0A86: rddata <= 8'h08;
            13'h0A87: rddata <= 8'hCD;
            13'h0A88: rddata <= 8'h37;
            13'h0A89: rddata <= 8'h0A;
            13'h0A8A: rddata <= 8'hE3;
            13'h0A8B: rddata <= 8'h11;
            13'h0A8C: rddata <= 8'h49;
            13'h0A8D: rddata <= 8'h0A;
            13'h0A8E: rddata <= 8'hD5;
            13'h0A8F: rddata <= 8'h01;
            13'h0A90: rddata <= 8'h15;
            13'h0A91: rddata <= 8'h02;
            13'h0A92: rddata <= 8'h09;
            13'h0A93: rddata <= 8'h4E;
            13'h0A94: rddata <= 8'h23;
            13'h0A95: rddata <= 8'h66;
            13'h0A96: rddata <= 8'h69;
            13'h0A97: rddata <= 8'hE9;
            13'h0A98: rddata <= 8'h15;
            13'h0A99: rddata <= 8'hFE;
            13'h0A9A: rddata <= 8'hA9;
            13'h0A9B: rddata <= 8'hC8;
            13'h0A9C: rddata <= 8'hFE;
            13'h0A9D: rddata <= 8'h2D;
            13'h0A9E: rddata <= 8'hC8;
            13'h0A9F: rddata <= 8'h14;
            13'h0AA0: rddata <= 8'hFE;
            13'h0AA1: rddata <= 8'h2B;
            13'h0AA2: rddata <= 8'hC8;
            13'h0AA3: rddata <= 8'hFE;
            13'h0AA4: rddata <= 8'hA8;
            13'h0AA5: rddata <= 8'hC8;
            13'h0AA6: rddata <= 8'h2B;
            13'h0AA7: rddata <= 8'hC9;
            13'h0AA8: rddata <= 8'hF6;
            13'h0AA9: rddata <= 8'hAF;
            13'h0AAA: rddata <= 8'hF5;
            13'h0AAB: rddata <= 8'hCD;
            13'h0AAC: rddata <= 8'h75;
            13'h0AAD: rddata <= 8'h09;
            13'h0AAE: rddata <= 8'hCD;
            13'h0AAF: rddata <= 8'h82;
            13'h0AB0: rddata <= 8'h06;
            13'h0AB1: rddata <= 8'hF1;
            13'h0AB2: rddata <= 8'hEB;
            13'h0AB3: rddata <= 8'hC1;
            13'h0AB4: rddata <= 8'hE3;
            13'h0AB5: rddata <= 8'hEB;
            13'h0AB6: rddata <= 8'hCD;
            13'h0AB7: rddata <= 8'h23;
            13'h0AB8: rddata <= 8'h15;
            13'h0AB9: rddata <= 8'hF5;
            13'h0ABA: rddata <= 8'hCD;
            13'h0ABB: rddata <= 8'h82;
            13'h0ABC: rddata <= 8'h06;
            13'h0ABD: rddata <= 8'hF1;
            13'h0ABE: rddata <= 8'hC1;
            13'h0ABF: rddata <= 8'h79;
            13'h0AC0: rddata <= 8'h21;
            13'h0AC1: rddata <= 8'h21;
            13'h0AC2: rddata <= 8'h0B;
            13'h0AC3: rddata <= 8'hC2;
            13'h0AC4: rddata <= 8'hCB;
            13'h0AC5: rddata <= 8'h0A;
            13'h0AC6: rddata <= 8'hA3;
            13'h0AC7: rddata <= 8'h4F;
            13'h0AC8: rddata <= 8'h78;
            13'h0AC9: rddata <= 8'hA2;
            13'h0ACA: rddata <= 8'hE9;
            13'h0ACB: rddata <= 8'hB3;
            13'h0ACC: rddata <= 8'h4F;
            13'h0ACD: rddata <= 8'h78;
            13'h0ACE: rddata <= 8'hB2;
            13'h0ACF: rddata <= 8'hE9;
            13'h0AD0: rddata <= 8'h21;
            13'h0AD1: rddata <= 8'hE2;
            13'h0AD2: rddata <= 8'h0A;
            13'h0AD3: rddata <= 8'h3A;
            13'h0AD4: rddata <= 8'hAB;
            13'h0AD5: rddata <= 8'h38;
            13'h0AD6: rddata <= 8'h1F;
            13'h0AD7: rddata <= 8'h7A;
            13'h0AD8: rddata <= 8'h17;
            13'h0AD9: rddata <= 8'h5F;
            13'h0ADA: rddata <= 8'h16;
            13'h0ADB: rddata <= 8'h64;
            13'h0ADC: rddata <= 8'h78;
            13'h0ADD: rddata <= 8'hBA;
            13'h0ADE: rddata <= 8'hD0;
            13'h0ADF: rddata <= 8'hC3;
            13'h0AE0: rddata <= 8'hCB;
            13'h0AE1: rddata <= 8'h09;
            13'h0AE2: rddata <= 8'hE4;
            13'h0AE3: rddata <= 8'h0A;
            13'h0AE4: rddata <= 8'h79;
            13'h0AE5: rddata <= 8'hB7;
            13'h0AE6: rddata <= 8'h1F;
            13'h0AE7: rddata <= 8'hC1;
            13'h0AE8: rddata <= 8'hD1;
            13'h0AE9: rddata <= 8'hF5;
            13'h0AEA: rddata <= 8'hCD;
            13'h0AEB: rddata <= 8'h77;
            13'h0AEC: rddata <= 8'h09;
            13'h0AED: rddata <= 8'h21;
            13'h0AEE: rddata <= 8'hFB;
            13'h0AEF: rddata <= 8'h0A;
            13'h0AF0: rddata <= 8'hE5;
            13'h0AF1: rddata <= 8'hCA;
            13'h0AF2: rddata <= 8'h5B;
            13'h0AF3: rddata <= 8'h15;
            13'h0AF4: rddata <= 8'hAF;
            13'h0AF5: rddata <= 8'h32;
            13'h0AF6: rddata <= 8'hAB;
            13'h0AF7: rddata <= 8'h38;
            13'h0AF8: rddata <= 8'hC3;
            13'h0AF9: rddata <= 8'hFC;
            13'h0AFA: rddata <= 8'h0D;
            13'h0AFB: rddata <= 8'h3C;
            13'h0AFC: rddata <= 8'h8F;
            13'h0AFD: rddata <= 8'hC1;
            13'h0AFE: rddata <= 8'hA0;
            13'h0AFF: rddata <= 8'hC6;
            13'h0B00: rddata <= 8'hFF;
            13'h0B01: rddata <= 8'h9F;
            13'h0B02: rddata <= 8'hC3;
            13'h0B03: rddata <= 8'hF6;
            13'h0B04: rddata <= 8'h14;
            13'h0B05: rddata <= 8'h16;
            13'h0B06: rddata <= 8'h5A;
            13'h0B07: rddata <= 8'hCD;
            13'h0B08: rddata <= 8'h88;
            13'h0B09: rddata <= 8'h09;
            13'h0B0A: rddata <= 8'hCD;
            13'h0B0B: rddata <= 8'h75;
            13'h0B0C: rddata <= 8'h09;
            13'h0B0D: rddata <= 8'hCD;
            13'h0B0E: rddata <= 8'h82;
            13'h0B0F: rddata <= 8'h06;
            13'h0B10: rddata <= 8'h7B;
            13'h0B11: rddata <= 8'h2F;
            13'h0B12: rddata <= 8'h4F;
            13'h0B13: rddata <= 8'h7A;
            13'h0B14: rddata <= 8'h2F;
            13'h0B15: rddata <= 8'hCD;
            13'h0B16: rddata <= 8'h21;
            13'h0B17: rddata <= 8'h0B;
            13'h0B18: rddata <= 8'hC1;
            13'h0B19: rddata <= 8'hC3;
            13'h0B1A: rddata <= 8'h94;
            13'h0B1B: rddata <= 8'h09;
            13'h0B1C: rddata <= 8'h7D;
            13'h0B1D: rddata <= 8'h93;
            13'h0B1E: rddata <= 8'h4F;
            13'h0B1F: rddata <= 8'h7C;
            13'h0B20: rddata <= 8'h9A;
            13'h0B21: rddata <= 8'h41;
            13'h0B22: rddata <= 8'h50;
            13'h0B23: rddata <= 8'h1E;
            13'h0B24: rddata <= 8'h00;
            13'h0B25: rddata <= 8'h21;
            13'h0B26: rddata <= 8'hAB;
            13'h0B27: rddata <= 8'h38;
            13'h0B28: rddata <= 8'h73;
            13'h0B29: rddata <= 8'h06;
            13'h0B2A: rddata <= 8'h90;
            13'h0B2B: rddata <= 8'hC3;
            13'h0B2C: rddata <= 8'hFB;
            13'h0B2D: rddata <= 8'h14;
            13'h0B2E: rddata <= 8'h3A;
            13'h0B2F: rddata <= 8'h46;
            13'h0B30: rddata <= 8'h38;
            13'h0B31: rddata <= 8'h18;
            13'h0B32: rddata <= 8'h03;
            13'h0B33: rddata <= 8'h3A;
            13'h0B34: rddata <= 8'h00;
            13'h0B35: rddata <= 8'h38;
            13'h0B36: rddata <= 8'h47;
            13'h0B37: rddata <= 8'hAF;
            13'h0B38: rddata <= 8'hC3;
            13'h0B39: rddata <= 8'h22;
            13'h0B3A: rddata <= 8'h0B;
            13'h0B3B: rddata <= 8'hF7;
            13'h0B3C: rddata <= 8'h0F;
            13'h0B3D: rddata <= 8'hC3;
            13'h0B3E: rddata <= 8'hC4;
            13'h0B3F: rddata <= 8'h03;
            13'h0B40: rddata <= 8'hF7;
            13'h0B41: rddata <= 8'h10;
            13'h0B42: rddata <= 8'hC3;
            13'h0B43: rddata <= 8'hC4;
            13'h0B44: rddata <= 8'h03;
            13'h0B45: rddata <= 8'hE5;
            13'h0B46: rddata <= 8'h2A;
            13'h0B47: rddata <= 8'h4D;
            13'h0B48: rddata <= 8'h38;
            13'h0B49: rddata <= 8'h23;
            13'h0B4A: rddata <= 8'h7C;
            13'h0B4B: rddata <= 8'hB5;
            13'h0B4C: rddata <= 8'hE1;
            13'h0B4D: rddata <= 8'hC0;
            13'h0B4E: rddata <= 8'h1E;
            13'h0B4F: rddata <= 8'h16;
            13'h0B50: rddata <= 8'hC3;
            13'h0B51: rddata <= 8'hDB;
            13'h0B52: rddata <= 8'h03;
            13'h0B53: rddata <= 8'hD7;
            13'h0B54: rddata <= 8'hCD;
            13'h0B55: rddata <= 8'h72;
            13'h0B56: rddata <= 8'h09;
            13'h0B57: rddata <= 8'hCD;
            13'h0B58: rddata <= 8'h7E;
            13'h0B59: rddata <= 8'h06;
            13'h0B5A: rddata <= 8'h7A;
            13'h0B5B: rddata <= 8'hB7;
            13'h0B5C: rddata <= 8'hC2;
            13'h0B5D: rddata <= 8'h97;
            13'h0B5E: rddata <= 8'h06;
            13'h0B5F: rddata <= 8'h2B;
            13'h0B60: rddata <= 8'hD7;
            13'h0B61: rddata <= 8'h7B;
            13'h0B62: rddata <= 8'hC9;
            13'h0B63: rddata <= 8'hCD;
            13'h0B64: rddata <= 8'h82;
            13'h0B65: rddata <= 8'h06;
            13'h0B66: rddata <= 8'hCD;
            13'h0B67: rddata <= 8'h88;
            13'h0B68: rddata <= 8'h0B;
            13'h0B69: rddata <= 8'h1A;
            13'h0B6A: rddata <= 8'hC3;
            13'h0B6B: rddata <= 8'h36;
            13'h0B6C: rddata <= 8'h0B;
            13'h0B6D: rddata <= 8'hCD;
            13'h0B6E: rddata <= 8'h72;
            13'h0B6F: rddata <= 8'h09;
            13'h0B70: rddata <= 8'hCD;
            13'h0B71: rddata <= 8'h82;
            13'h0B72: rddata <= 8'h06;
            13'h0B73: rddata <= 8'hCD;
            13'h0B74: rddata <= 8'h88;
            13'h0B75: rddata <= 8'h0B;
            13'h0B76: rddata <= 8'hD5;
            13'h0B77: rddata <= 8'hCF;
            13'h0B78: rddata <= 8'h2C;
            13'h0B79: rddata <= 8'hCD;
            13'h0B7A: rddata <= 8'h54;
            13'h0B7B: rddata <= 8'h0B;
            13'h0B7C: rddata <= 8'hD1;
            13'h0B7D: rddata <= 8'h12;
            13'h0B7E: rddata <= 8'hC9;
            13'h0B7F: rddata <= 8'hCD;
            13'h0B80: rddata <= 8'h85;
            13'h0B81: rddata <= 8'h09;
            13'h0B82: rddata <= 8'hE5;
            13'h0B83: rddata <= 8'hCD;
            13'h0B84: rddata <= 8'h82;
            13'h0B85: rddata <= 8'h06;
            13'h0B86: rddata <= 8'hE1;
            13'h0B87: rddata <= 8'hC9;
            13'h0B88: rddata <= 8'hE5;
            13'h0B89: rddata <= 8'h21;
            13'h0B8A: rddata <= 8'hFF;
            13'h0B8B: rddata <= 8'h2F;
            13'h0B8C: rddata <= 8'hE7;
            13'h0B8D: rddata <= 8'hE1;
            13'h0B8E: rddata <= 8'hD2;
            13'h0B8F: rddata <= 8'h97;
            13'h0B90: rddata <= 8'h06;
            13'h0B91: rddata <= 8'hC9;
            13'h0B92: rddata <= 8'hCD;
            13'h0B93: rddata <= 8'hA9;
            13'h0B94: rddata <= 8'h0B;
            13'h0B95: rddata <= 8'hC5;
            13'h0B96: rddata <= 8'hE3;
            13'h0B97: rddata <= 8'hC1;
            13'h0B98: rddata <= 8'hE7;
            13'h0B99: rddata <= 8'h7E;
            13'h0B9A: rddata <= 8'h02;
            13'h0B9B: rddata <= 8'hC8;
            13'h0B9C: rddata <= 8'h0B;
            13'h0B9D: rddata <= 8'h2B;
            13'h0B9E: rddata <= 8'h18;
            13'h0B9F: rddata <= 8'hF8;
            13'h0BA0: rddata <= 8'hE5;
            13'h0BA1: rddata <= 8'h2A;
            13'h0BA2: rddata <= 8'hDA;
            13'h0BA3: rddata <= 8'h38;
            13'h0BA4: rddata <= 8'h06;
            13'h0BA5: rddata <= 8'h00;
            13'h0BA6: rddata <= 8'h09;
            13'h0BA7: rddata <= 8'h09;
            13'h0BA8: rddata <= 8'h3E;
            13'h0BA9: rddata <= 8'hE5;
            13'h0BAA: rddata <= 8'h3E;
            13'h0BAB: rddata <= 8'hD0;
            13'h0BAC: rddata <= 8'h95;
            13'h0BAD: rddata <= 8'h6F;
            13'h0BAE: rddata <= 8'h3E;
            13'h0BAF: rddata <= 8'hFF;
            13'h0BB0: rddata <= 8'h9C;
            13'h0BB1: rddata <= 8'h67;
            13'h0BB2: rddata <= 8'h38;
            13'h0BB3: rddata <= 8'h03;
            13'h0BB4: rddata <= 8'h39;
            13'h0BB5: rddata <= 8'hE1;
            13'h0BB6: rddata <= 8'hD8;
            13'h0BB7: rddata <= 8'h11;
            13'h0BB8: rddata <= 8'h0C;
            13'h0BB9: rddata <= 8'h00;
            13'h0BBA: rddata <= 8'hC3;
            13'h0BBB: rddata <= 8'hDB;
            13'h0BBC: rddata <= 8'h03;
            13'h0BBD: rddata <= 8'hC0;
            13'h0BBE: rddata <= 8'hF7;
            13'h0BBF: rddata <= 8'h0C;
            13'h0BC0: rddata <= 8'h2A;
            13'h0BC1: rddata <= 8'h4F;
            13'h0BC2: rddata <= 8'h38;
            13'h0BC3: rddata <= 8'hAF;
            13'h0BC4: rddata <= 8'h77;
            13'h0BC5: rddata <= 8'h23;
            13'h0BC6: rddata <= 8'h77;
            13'h0BC7: rddata <= 8'h23;
            13'h0BC8: rddata <= 8'h22;
            13'h0BC9: rddata <= 8'hD6;
            13'h0BCA: rddata <= 8'h38;
            13'h0BCB: rddata <= 8'h2A;
            13'h0BCC: rddata <= 8'h4F;
            13'h0BCD: rddata <= 8'h38;
            13'h0BCE: rddata <= 8'h2B;
            13'h0BCF: rddata <= 8'h22;
            13'h0BD0: rddata <= 8'hCE;
            13'h0BD1: rddata <= 8'h38;
            13'h0BD2: rddata <= 8'h2A;
            13'h0BD3: rddata <= 8'hAD;
            13'h0BD4: rddata <= 8'h38;
            13'h0BD5: rddata <= 8'h22;
            13'h0BD6: rddata <= 8'hC1;
            13'h0BD7: rddata <= 8'h38;
            13'h0BD8: rddata <= 8'hAF;
            13'h0BD9: rddata <= 8'hCD;
            13'h0BDA: rddata <= 8'h05;
            13'h0BDB: rddata <= 8'h0C;
            13'h0BDC: rddata <= 8'h2A;
            13'h0BDD: rddata <= 8'hD6;
            13'h0BDE: rddata <= 8'h38;
            13'h0BDF: rddata <= 8'h22;
            13'h0BE0: rddata <= 8'hD8;
            13'h0BE1: rddata <= 8'h38;
            13'h0BE2: rddata <= 8'h22;
            13'h0BE3: rddata <= 8'hDA;
            13'h0BE4: rddata <= 8'h38;
            13'h0BE5: rddata <= 8'hC1;
            13'h0BE6: rddata <= 8'h2A;
            13'h0BE7: rddata <= 8'h4B;
            13'h0BE8: rddata <= 8'h38;
            13'h0BE9: rddata <= 8'hF9;
            13'h0BEA: rddata <= 8'hCD;
            13'h0BEB: rddata <= 8'hD8;
            13'h0BEC: rddata <= 8'h1F;
            13'h0BED: rddata <= 8'h22;
            13'h0BEE: rddata <= 8'hAF;
            13'h0BEF: rddata <= 8'h38;
            13'h0BF0: rddata <= 8'hCD;
            13'h0BF1: rddata <= 8'hBE;
            13'h0BF2: rddata <= 8'h19;
            13'h0BF3: rddata <= 8'hAF;
            13'h0BF4: rddata <= 8'h6F;
            13'h0BF5: rddata <= 8'h67;
            13'h0BF6: rddata <= 8'h22;
            13'h0BF7: rddata <= 8'hD4;
            13'h0BF8: rddata <= 8'h38;
            13'h0BF9: rddata <= 8'h32;
            13'h0BFA: rddata <= 8'hCB;
            13'h0BFB: rddata <= 8'h38;
            13'h0BFC: rddata <= 8'h22;
            13'h0BFD: rddata <= 8'hDE;
            13'h0BFE: rddata <= 8'h38;
            13'h0BFF: rddata <= 8'hE5;
            13'h0C00: rddata <= 8'hC5;
            13'h0C01: rddata <= 8'h2A;
            13'h0C02: rddata <= 8'hCE;
            13'h0C03: rddata <= 8'h38;
            13'h0C04: rddata <= 8'hC9;
            13'h0C05: rddata <= 8'hEB;
            13'h0C06: rddata <= 8'h2A;
            13'h0C07: rddata <= 8'h4F;
            13'h0C08: rddata <= 8'h38;
            13'h0C09: rddata <= 8'h28;
            13'h0C0A: rddata <= 8'h0E;
            13'h0C0B: rddata <= 8'hEB;
            13'h0C0C: rddata <= 8'hCD;
            13'h0C0D: rddata <= 8'h9C;
            13'h0C0E: rddata <= 8'h06;
            13'h0C0F: rddata <= 8'hE5;
            13'h0C10: rddata <= 8'hCD;
            13'h0C11: rddata <= 8'h9F;
            13'h0C12: rddata <= 8'h04;
            13'h0C13: rddata <= 8'h60;
            13'h0C14: rddata <= 8'h69;
            13'h0C15: rddata <= 8'hD1;
            13'h0C16: rddata <= 8'hD2;
            13'h0C17: rddata <= 8'hF3;
            13'h0C18: rddata <= 8'h06;
            13'h0C19: rddata <= 8'h2B;
            13'h0C1A: rddata <= 8'h22;
            13'h0C1B: rddata <= 8'hDC;
            13'h0C1C: rddata <= 8'h38;
            13'h0C1D: rddata <= 8'hEB;
            13'h0C1E: rddata <= 8'hC9;
            13'h0C1F: rddata <= 8'hC0;
            13'h0C20: rddata <= 8'hF6;
            13'h0C21: rddata <= 8'hC0;
            13'h0C22: rddata <= 8'h22;
            13'h0C23: rddata <= 8'hCE;
            13'h0C24: rddata <= 8'h38;
            13'h0C25: rddata <= 8'h21;
            13'h0C26: rddata <= 8'hF6;
            13'h0C27: rddata <= 8'hFF;
            13'h0C28: rddata <= 8'hC1;
            13'h0C29: rddata <= 8'h2A;
            13'h0C2A: rddata <= 8'h4D;
            13'h0C2B: rddata <= 8'h38;
            13'h0C2C: rddata <= 8'hF5;
            13'h0C2D: rddata <= 8'h7D;
            13'h0C2E: rddata <= 8'hA4;
            13'h0C2F: rddata <= 8'h3C;
            13'h0C30: rddata <= 8'h28;
            13'h0C31: rddata <= 8'h09;
            13'h0C32: rddata <= 8'h22;
            13'h0C33: rddata <= 8'hD2;
            13'h0C34: rddata <= 8'h38;
            13'h0C35: rddata <= 8'h2A;
            13'h0C36: rddata <= 8'hCE;
            13'h0C37: rddata <= 8'h38;
            13'h0C38: rddata <= 8'h22;
            13'h0C39: rddata <= 8'hD4;
            13'h0C3A: rddata <= 8'h38;
            13'h0C3B: rddata <= 8'hCD;
            13'h0C3C: rddata <= 8'hBE;
            13'h0C3D: rddata <= 8'h19;
            13'h0C3E: rddata <= 8'hCD;
            13'h0C3F: rddata <= 8'hDE;
            13'h0C40: rddata <= 8'h19;
            13'h0C41: rddata <= 8'hF1;
            13'h0C42: rddata <= 8'h21;
            13'h0C43: rddata <= 8'h73;
            13'h0C44: rddata <= 8'h03;
            13'h0C45: rddata <= 8'hC2;
            13'h0C46: rddata <= 8'hF4;
            13'h0C47: rddata <= 8'h03;
            13'h0C48: rddata <= 8'hC3;
            13'h0C49: rddata <= 8'h02;
            13'h0C4A: rddata <= 8'h04;
            13'h0C4B: rddata <= 8'h2A;
            13'h0C4C: rddata <= 8'hD4;
            13'h0C4D: rddata <= 8'h38;
            13'h0C4E: rddata <= 8'h7C;
            13'h0C4F: rddata <= 8'hB5;
            13'h0C50: rddata <= 8'h11;
            13'h0C51: rddata <= 8'h20;
            13'h0C52: rddata <= 8'h00;
            13'h0C53: rddata <= 8'hCA;
            13'h0C54: rddata <= 8'hDB;
            13'h0C55: rddata <= 8'h03;
            13'h0C56: rddata <= 8'hED;
            13'h0C57: rddata <= 8'h5B;
            13'h0C58: rddata <= 8'hD2;
            13'h0C59: rddata <= 8'h38;
            13'h0C5A: rddata <= 8'hED;
            13'h0C5B: rddata <= 8'h53;
            13'h0C5C: rddata <= 8'h4D;
            13'h0C5D: rddata <= 8'h38;
            13'h0C5E: rddata <= 8'hC9;
            13'h0C5F: rddata <= 8'hC3;
            13'h0C60: rddata <= 8'h97;
            13'h0C61: rddata <= 8'h06;
            13'h0C62: rddata <= 8'h3E;
            13'h0C63: rddata <= 8'hAF;
            13'h0C64: rddata <= 8'hB7;
            13'h0C65: rddata <= 8'hF5;
            13'h0C66: rddata <= 8'hD7;
            13'h0C67: rddata <= 8'h3E;
            13'h0C68: rddata <= 8'h01;
            13'h0C69: rddata <= 8'h32;
            13'h0C6A: rddata <= 8'hCB;
            13'h0C6B: rddata <= 8'h38;
            13'h0C6C: rddata <= 8'hCD;
            13'h0C6D: rddata <= 8'hD1;
            13'h0C6E: rddata <= 8'h10;
            13'h0C6F: rddata <= 8'hC2;
            13'h0C70: rddata <= 8'h97;
            13'h0C71: rddata <= 8'h06;
            13'h0C72: rddata <= 8'h32;
            13'h0C73: rddata <= 8'hCB;
            13'h0C74: rddata <= 8'h38;
            13'h0C75: rddata <= 8'hCD;
            13'h0C76: rddata <= 8'h75;
            13'h0C77: rddata <= 8'h09;
            13'h0C78: rddata <= 8'hF1;
            13'h0C79: rddata <= 8'hE5;
            13'h0C7A: rddata <= 8'hF5;
            13'h0C7B: rddata <= 8'hC5;
            13'h0C7C: rddata <= 8'h06;
            13'h0C7D: rddata <= 8'h23;
            13'h0C7E: rddata <= 8'h28;
            13'h0C7F: rddata <= 8'h12;
            13'h0C80: rddata <= 8'hCD;
            13'h0C81: rddata <= 8'h7F;
            13'h0C82: rddata <= 8'h1B;
            13'h0C83: rddata <= 8'hCD;
            13'h0C84: rddata <= 8'hBC;
            13'h0C85: rddata <= 8'h1B;
            13'h0C86: rddata <= 8'h78;
            13'h0C87: rddata <= 8'hCD;
            13'h0C88: rddata <= 8'h87;
            13'h0C89: rddata <= 8'h1B;
            13'h0C8A: rddata <= 8'hCD;
            13'h0C8B: rddata <= 8'h87;
            13'h0C8C: rddata <= 8'h1B;
            13'h0C8D: rddata <= 8'hCD;
            13'h0C8E: rddata <= 8'h87;
            13'h0C8F: rddata <= 8'h1B;
            13'h0C90: rddata <= 8'h18;
            13'h0C91: rddata <= 8'h11;
            13'h0C92: rddata <= 8'hCD;
            13'h0C93: rddata <= 8'h2E;
            13'h0C94: rddata <= 8'h1B;
            13'h0C95: rddata <= 8'hCD;
            13'h0C96: rddata <= 8'hCE;
            13'h0C97: rddata <= 8'h1B;
            13'h0C98: rddata <= 8'h0E;
            13'h0C99: rddata <= 8'h06;
            13'h0C9A: rddata <= 8'hCD;
            13'h0C9B: rddata <= 8'h4D;
            13'h0C9C: rddata <= 8'h1B;
            13'h0C9D: rddata <= 8'hB8;
            13'h0C9E: rddata <= 8'h20;
            13'h0C9F: rddata <= 8'hF8;
            13'h0CA0: rddata <= 8'h0D;
            13'h0CA1: rddata <= 8'h20;
            13'h0CA2: rddata <= 8'hF7;
            13'h0CA3: rddata <= 8'hE1;
            13'h0CA4: rddata <= 8'hEB;
            13'h0CA5: rddata <= 8'h19;
            13'h0CA6: rddata <= 8'hEB;
            13'h0CA7: rddata <= 8'h4E;
            13'h0CA8: rddata <= 8'h06;
            13'h0CA9: rddata <= 8'h00;
            13'h0CAA: rddata <= 8'h09;
            13'h0CAB: rddata <= 8'h09;
            13'h0CAC: rddata <= 8'h23;
            13'h0CAD: rddata <= 8'hE7;
            13'h0CAE: rddata <= 8'h28;
            13'h0CAF: rddata <= 8'h0D;
            13'h0CB0: rddata <= 8'hF1;
            13'h0CB1: rddata <= 8'hF5;
            13'h0CB2: rddata <= 8'h7E;
            13'h0CB3: rddata <= 8'hC4;
            13'h0CB4: rddata <= 8'h8A;
            13'h0CB5: rddata <= 8'h1B;
            13'h0CB6: rddata <= 8'hCC;
            13'h0CB7: rddata <= 8'h4D;
            13'h0CB8: rddata <= 8'h1B;
            13'h0CB9: rddata <= 8'h77;
            13'h0CBA: rddata <= 8'h23;
            13'h0CBB: rddata <= 8'h18;
            13'h0CBC: rddata <= 8'hF0;
            13'h0CBD: rddata <= 8'hF1;
            13'h0CBE: rddata <= 8'hC2;
            13'h0CBF: rddata <= 8'h1C;
            13'h0CC0: rddata <= 8'h1C;
            13'h0CC1: rddata <= 8'hE1;
            13'h0CC2: rddata <= 8'hC3;
            13'h0CC3: rddata <= 8'h7E;
            13'h0CC4: rddata <= 8'h1B;
            13'h0CC5: rddata <= 8'h7E;
            13'h0CC6: rddata <= 8'hFE;
            13'h0CC7: rddata <= 8'h41;
            13'h0CC8: rddata <= 8'hD8;
            13'h0CC9: rddata <= 8'hFE;
            13'h0CCA: rddata <= 8'h5B;
            13'h0CCB: rddata <= 8'h3F;
            13'h0CCC: rddata <= 8'hC9;
            13'h0CCD: rddata <= 8'hF7;
            13'h0CCE: rddata <= 8'h0B;
            13'h0CCF: rddata <= 8'hCA;
            13'h0CD0: rddata <= 8'hCF;
            13'h0CD1: rddata <= 8'h0B;
            13'h0CD2: rddata <= 8'hCD;
            13'h0CD3: rddata <= 8'h7B;
            13'h0CD4: rddata <= 8'h06;
            13'h0CD5: rddata <= 8'h2B;
            13'h0CD6: rddata <= 8'hD7;
            13'h0CD7: rddata <= 8'hE5;
            13'h0CD8: rddata <= 8'h2A;
            13'h0CD9: rddata <= 8'hAD;
            13'h0CDA: rddata <= 8'h38;
            13'h0CDB: rddata <= 8'h28;
            13'h0CDC: rddata <= 8'h0E;
            13'h0CDD: rddata <= 8'hE1;
            13'h0CDE: rddata <= 8'hCF;
            13'h0CDF: rddata <= 8'h2C;
            13'h0CE0: rddata <= 8'hD5;
            13'h0CE1: rddata <= 8'hCD;
            13'h0CE2: rddata <= 8'h7B;
            13'h0CE3: rddata <= 8'h06;
            13'h0CE4: rddata <= 8'h2B;
            13'h0CE5: rddata <= 8'hD7;
            13'h0CE6: rddata <= 8'hC2;
            13'h0CE7: rddata <= 8'hC4;
            13'h0CE8: rddata <= 8'h03;
            13'h0CE9: rddata <= 8'hE3;
            13'h0CEA: rddata <= 8'hEB;
            13'h0CEB: rddata <= 8'h7D;
            13'h0CEC: rddata <= 8'h93;
            13'h0CED: rddata <= 8'h5F;
            13'h0CEE: rddata <= 8'h7C;
            13'h0CEF: rddata <= 8'h9A;
            13'h0CF0: rddata <= 8'h57;
            13'h0CF1: rddata <= 8'hDA;
            13'h0CF2: rddata <= 8'hB7;
            13'h0CF3: rddata <= 8'h0B;
            13'h0CF4: rddata <= 8'hE5;
            13'h0CF5: rddata <= 8'h2A;
            13'h0CF6: rddata <= 8'hD6;
            13'h0CF7: rddata <= 8'h38;
            13'h0CF8: rddata <= 8'h01;
            13'h0CF9: rddata <= 8'h28;
            13'h0CFA: rddata <= 8'h00;
            13'h0CFB: rddata <= 8'h09;
            13'h0CFC: rddata <= 8'hE7;
            13'h0CFD: rddata <= 8'hD2;
            13'h0CFE: rddata <= 8'hB7;
            13'h0CFF: rddata <= 8'h0B;
            13'h0D00: rddata <= 8'hEB;
            13'h0D01: rddata <= 8'h22;
            13'h0D02: rddata <= 8'h4B;
            13'h0D03: rddata <= 8'h38;
            13'h0D04: rddata <= 8'hE1;
            13'h0D05: rddata <= 8'h22;
            13'h0D06: rddata <= 8'hAD;
            13'h0D07: rddata <= 8'h38;
            13'h0D08: rddata <= 8'hE1;
            13'h0D09: rddata <= 8'hC3;
            13'h0D0A: rddata <= 8'hCF;
            13'h0D0B: rddata <= 8'h0B;
            13'h0D0C: rddata <= 8'h7D;
            13'h0D0D: rddata <= 8'h93;
            13'h0D0E: rddata <= 8'h5F;
            13'h0D0F: rddata <= 8'h7C;
            13'h0D10: rddata <= 8'h9A;
            13'h0D11: rddata <= 8'h57;
            13'h0D12: rddata <= 8'hC9;
            13'h0D13: rddata <= 8'h11;
            13'h0D14: rddata <= 8'h00;
            13'h0D15: rddata <= 8'h00;
            13'h0D16: rddata <= 8'hC4;
            13'h0D17: rddata <= 8'hD1;
            13'h0D18: rddata <= 8'h10;
            13'h0D19: rddata <= 8'h22;
            13'h0D1A: rddata <= 8'hCE;
            13'h0D1B: rddata <= 8'h38;
            13'h0D1C: rddata <= 8'hCD;
            13'h0D1D: rddata <= 8'h9F;
            13'h0D1E: rddata <= 8'h03;
            13'h0D1F: rddata <= 8'hC2;
            13'h0D20: rddata <= 8'hCA;
            13'h0D21: rddata <= 8'h03;
            13'h0D22: rddata <= 8'hF9;
            13'h0D23: rddata <= 8'hD5;
            13'h0D24: rddata <= 8'h7E;
            13'h0D25: rddata <= 8'hF5;
            13'h0D26: rddata <= 8'h23;
            13'h0D27: rddata <= 8'hD5;
            13'h0D28: rddata <= 8'hCD;
            13'h0D29: rddata <= 8'h20;
            13'h0D2A: rddata <= 8'h15;
            13'h0D2B: rddata <= 8'hE3;
            13'h0D2C: rddata <= 8'hE5;
            13'h0D2D: rddata <= 8'hCD;
            13'h0D2E: rddata <= 8'h53;
            13'h0D2F: rddata <= 8'h12;
            13'h0D30: rddata <= 8'hE1;
            13'h0D31: rddata <= 8'hCD;
            13'h0D32: rddata <= 8'h3A;
            13'h0D33: rddata <= 8'h15;
            13'h0D34: rddata <= 8'hE1;
            13'h0D35: rddata <= 8'hCD;
            13'h0D36: rddata <= 8'h31;
            13'h0D37: rddata <= 8'h15;
            13'h0D38: rddata <= 8'hE5;
            13'h0D39: rddata <= 8'hCD;
            13'h0D3A: rddata <= 8'h5B;
            13'h0D3B: rddata <= 8'h15;
            13'h0D3C: rddata <= 8'hE1;
            13'h0D3D: rddata <= 8'hC1;
            13'h0D3E: rddata <= 8'h90;
            13'h0D3F: rddata <= 8'hCD;
            13'h0D40: rddata <= 8'h31;
            13'h0D41: rddata <= 8'h15;
            13'h0D42: rddata <= 8'h28;
            13'h0D43: rddata <= 8'h09;
            13'h0D44: rddata <= 8'hEB;
            13'h0D45: rddata <= 8'h22;
            13'h0D46: rddata <= 8'h4D;
            13'h0D47: rddata <= 8'h38;
            13'h0D48: rddata <= 8'h69;
            13'h0D49: rddata <= 8'h60;
            13'h0D4A: rddata <= 8'hC3;
            13'h0D4B: rddata <= 8'h28;
            13'h0D4C: rddata <= 8'h06;
            13'h0D4D: rddata <= 8'hF9;
            13'h0D4E: rddata <= 8'h2A;
            13'h0D4F: rddata <= 8'hCE;
            13'h0D50: rddata <= 8'h38;
            13'h0D51: rddata <= 8'h7E;
            13'h0D52: rddata <= 8'hFE;
            13'h0D53: rddata <= 8'h2C;
            13'h0D54: rddata <= 8'hC2;
            13'h0D55: rddata <= 8'h2C;
            13'h0D56: rddata <= 8'h06;
            13'h0D57: rddata <= 8'hD7;
            13'h0D58: rddata <= 8'hCD;
            13'h0D59: rddata <= 8'h16;
            13'h0D5A: rddata <= 8'h0D;
            13'h0D5B: rddata <= 8'h3E;
            13'h0D5C: rddata <= 8'h3F;
            13'h0D5D: rddata <= 8'hDF;
            13'h0D5E: rddata <= 8'h3E;
            13'h0D5F: rddata <= 8'h20;
            13'h0D60: rddata <= 8'hDF;
            13'h0D61: rddata <= 8'hC3;
            13'h0D62: rddata <= 8'h85;
            13'h0D63: rddata <= 8'h0D;
            13'h0D64: rddata <= 8'h3A;
            13'h0D65: rddata <= 8'h4A;
            13'h0D66: rddata <= 8'h38;
            13'h0D67: rddata <= 8'hB7;
            13'h0D68: rddata <= 8'h3E;
            13'h0D69: rddata <= 8'h5C;
            13'h0D6A: rddata <= 8'h32;
            13'h0D6B: rddata <= 8'h4A;
            13'h0D6C: rddata <= 8'h38;
            13'h0D6D: rddata <= 8'h20;
            13'h0D6E: rddata <= 8'h05;
            13'h0D6F: rddata <= 8'h05;
            13'h0D70: rddata <= 8'h28;
            13'h0D71: rddata <= 8'h13;
            13'h0D72: rddata <= 8'hDF;
            13'h0D73: rddata <= 8'h04;
            13'h0D74: rddata <= 8'h05;
            13'h0D75: rddata <= 8'h2B;
            13'h0D76: rddata <= 8'h28;
            13'h0D77: rddata <= 8'h09;
            13'h0D78: rddata <= 8'h7E;
            13'h0D79: rddata <= 8'hDF;
            13'h0D7A: rddata <= 8'h18;
            13'h0D7B: rddata <= 8'h12;
            13'h0D7C: rddata <= 8'h05;
            13'h0D7D: rddata <= 8'h2B;
            13'h0D7E: rddata <= 8'hDF;
            13'h0D7F: rddata <= 8'h20;
            13'h0D80: rddata <= 8'h0D;
            13'h0D81: rddata <= 8'hDF;
            13'h0D82: rddata <= 8'hCD;
            13'h0D83: rddata <= 8'hEA;
            13'h0D84: rddata <= 8'h19;
            13'h0D85: rddata <= 8'h21;
            13'h0D86: rddata <= 8'h60;
            13'h0D87: rddata <= 8'h38;
            13'h0D88: rddata <= 8'h06;
            13'h0D89: rddata <= 8'h01;
            13'h0D8A: rddata <= 8'hAF;
            13'h0D8B: rddata <= 8'h32;
            13'h0D8C: rddata <= 8'h4A;
            13'h0D8D: rddata <= 8'h38;
            13'h0D8E: rddata <= 8'hCD;
            13'h0D8F: rddata <= 8'hDA;
            13'h0D90: rddata <= 8'h19;
            13'h0D91: rddata <= 8'h4F;
            13'h0D92: rddata <= 8'hFE;
            13'h0D93: rddata <= 8'h7F;
            13'h0D94: rddata <= 8'h28;
            13'h0D95: rddata <= 8'hCE;
            13'h0D96: rddata <= 8'h3A;
            13'h0D97: rddata <= 8'h4A;
            13'h0D98: rddata <= 8'h38;
            13'h0D99: rddata <= 8'hB7;
            13'h0D9A: rddata <= 8'h28;
            13'h0D9B: rddata <= 8'h07;
            13'h0D9C: rddata <= 8'h3E;
            13'h0D9D: rddata <= 8'h5C;
            13'h0D9E: rddata <= 8'hDF;
            13'h0D9F: rddata <= 8'hAF;
            13'h0DA0: rddata <= 8'h32;
            13'h0DA1: rddata <= 8'h4A;
            13'h0DA2: rddata <= 8'h38;
            13'h0DA3: rddata <= 8'h79;
            13'h0DA4: rddata <= 8'hFE;
            13'h0DA5: rddata <= 8'h07;
            13'h0DA6: rddata <= 8'h28;
            13'h0DA7: rddata <= 8'h41;
            13'h0DA8: rddata <= 8'hFE;
            13'h0DA9: rddata <= 8'h03;
            13'h0DAA: rddata <= 8'hCC;
            13'h0DAB: rddata <= 8'hEA;
            13'h0DAC: rddata <= 8'h19;
            13'h0DAD: rddata <= 8'h37;
            13'h0DAE: rddata <= 8'hC8;
            13'h0DAF: rddata <= 8'hFE;
            13'h0DB0: rddata <= 8'h0D;
            13'h0DB1: rddata <= 8'hCA;
            13'h0DB2: rddata <= 8'hE5;
            13'h0DB3: rddata <= 8'h19;
            13'h0DB4: rddata <= 8'hFE;
            13'h0DB5: rddata <= 8'h15;
            13'h0DB6: rddata <= 8'hCA;
            13'h0DB7: rddata <= 8'h82;
            13'h0DB8: rddata <= 8'h0D;
            13'h0DB9: rddata <= 8'h00;
            13'h0DBA: rddata <= 8'h00;
            13'h0DBB: rddata <= 8'h00;
            13'h0DBC: rddata <= 8'h00;
            13'h0DBD: rddata <= 8'h00;
            13'h0DBE: rddata <= 8'hFE;
            13'h0DBF: rddata <= 8'h08;
            13'h0DC0: rddata <= 8'hCA;
            13'h0DC1: rddata <= 8'h7C;
            13'h0DC2: rddata <= 8'h0D;
            13'h0DC3: rddata <= 8'hFE;
            13'h0DC4: rddata <= 8'h18;
            13'h0DC5: rddata <= 8'h20;
            13'h0DC6: rddata <= 8'h05;
            13'h0DC7: rddata <= 8'h3E;
            13'h0DC8: rddata <= 8'h23;
            13'h0DC9: rddata <= 8'hC3;
            13'h0DCA: rddata <= 8'h81;
            13'h0DCB: rddata <= 8'h0D;
            13'h0DCC: rddata <= 8'hFE;
            13'h0DCD: rddata <= 8'h12;
            13'h0DCE: rddata <= 8'h20;
            13'h0DCF: rddata <= 8'h14;
            13'h0DD0: rddata <= 8'hC5;
            13'h0DD1: rddata <= 8'hD5;
            13'h0DD2: rddata <= 8'hE5;
            13'h0DD3: rddata <= 8'h36;
            13'h0DD4: rddata <= 8'h00;
            13'h0DD5: rddata <= 8'hCD;
            13'h0DD6: rddata <= 8'hEA;
            13'h0DD7: rddata <= 8'h19;
            13'h0DD8: rddata <= 8'h21;
            13'h0DD9: rddata <= 8'h60;
            13'h0DDA: rddata <= 8'h38;
            13'h0DDB: rddata <= 8'hCD;
            13'h0DDC: rddata <= 8'h9D;
            13'h0DDD: rddata <= 8'h0E;
            13'h0DDE: rddata <= 8'hE1;
            13'h0DDF: rddata <= 8'hD1;
            13'h0DE0: rddata <= 8'hC1;
            13'h0DE1: rddata <= 8'hC3;
            13'h0DE2: rddata <= 8'h8E;
            13'h0DE3: rddata <= 8'h0D;
            13'h0DE4: rddata <= 8'hFE;
            13'h0DE5: rddata <= 8'h20;
            13'h0DE6: rddata <= 8'hDA;
            13'h0DE7: rddata <= 8'h8E;
            13'h0DE8: rddata <= 8'h0D;
            13'h0DE9: rddata <= 8'h78;
            13'h0DEA: rddata <= 8'hFE;
            13'h0DEB: rddata <= 8'h49;
            13'h0DEC: rddata <= 8'h3E;
            13'h0DED: rddata <= 8'h07;
            13'h0DEE: rddata <= 8'hD2;
            13'h0DEF: rddata <= 8'hF8;
            13'h0DF0: rddata <= 8'h0D;
            13'h0DF1: rddata <= 8'h79;
            13'h0DF2: rddata <= 8'h71;
            13'h0DF3: rddata <= 8'h32;
            13'h0DF4: rddata <= 8'hCC;
            13'h0DF5: rddata <= 8'h38;
            13'h0DF6: rddata <= 8'h23;
            13'h0DF7: rddata <= 8'h04;
            13'h0DF8: rddata <= 8'hDF;
            13'h0DF9: rddata <= 8'hC3;
            13'h0DFA: rddata <= 8'h8E;
            13'h0DFB: rddata <= 8'h0D;
            13'h0DFC: rddata <= 8'hD5;
            13'h0DFD: rddata <= 8'hCD;
            13'h0DFE: rddata <= 8'hC9;
            13'h0DFF: rddata <= 8'h0F;
            13'h0E00: rddata <= 8'h7E;
            13'h0E01: rddata <= 8'h23;
            13'h0E02: rddata <= 8'h23;
            13'h0E03: rddata <= 8'h4E;
            13'h0E04: rddata <= 8'h23;
            13'h0E05: rddata <= 8'h46;
            13'h0E06: rddata <= 8'hD1;
            13'h0E07: rddata <= 8'hC5;
            13'h0E08: rddata <= 8'hF5;
            13'h0E09: rddata <= 8'hCD;
            13'h0E0A: rddata <= 8'hCD;
            13'h0E0B: rddata <= 8'h0F;
            13'h0E0C: rddata <= 8'hCD;
            13'h0E0D: rddata <= 8'h31;
            13'h0E0E: rddata <= 8'h15;
            13'h0E0F: rddata <= 8'hF1;
            13'h0E10: rddata <= 8'h57;
            13'h0E11: rddata <= 8'hE1;
            13'h0E12: rddata <= 8'h7B;
            13'h0E13: rddata <= 8'hB2;
            13'h0E14: rddata <= 8'hC8;
            13'h0E15: rddata <= 8'h7A;
            13'h0E16: rddata <= 8'hD6;
            13'h0E17: rddata <= 8'h01;
            13'h0E18: rddata <= 8'hD8;
            13'h0E19: rddata <= 8'hAF;
            13'h0E1A: rddata <= 8'hBB;
            13'h0E1B: rddata <= 8'h3C;
            13'h0E1C: rddata <= 8'hD0;
            13'h0E1D: rddata <= 8'h15;
            13'h0E1E: rddata <= 8'h1D;
            13'h0E1F: rddata <= 8'h0A;
            13'h0E20: rddata <= 8'h03;
            13'h0E21: rddata <= 8'hBE;
            13'h0E22: rddata <= 8'h23;
            13'h0E23: rddata <= 8'h28;
            13'h0E24: rddata <= 8'hED;
            13'h0E25: rddata <= 8'h3F;
            13'h0E26: rddata <= 8'hC3;
            13'h0E27: rddata <= 8'hF1;
            13'h0E28: rddata <= 8'h14;
            13'h0E29: rddata <= 8'hCD;
            13'h0E2A: rddata <= 8'h75;
            13'h0E2B: rddata <= 8'h09;
            13'h0E2C: rddata <= 8'hCD;
            13'h0E2D: rddata <= 8'h80;
            13'h0E2E: rddata <= 8'h16;
            13'h0E2F: rddata <= 8'hCD;
            13'h0E30: rddata <= 8'h5F;
            13'h0E31: rddata <= 8'h0E;
            13'h0E32: rddata <= 8'hCD;
            13'h0E33: rddata <= 8'hC9;
            13'h0E34: rddata <= 8'h0F;
            13'h0E35: rddata <= 8'h01;
            13'h0E36: rddata <= 8'h1D;
            13'h0E37: rddata <= 8'h10;
            13'h0E38: rddata <= 8'hC5;
            13'h0E39: rddata <= 8'h7E;
            13'h0E3A: rddata <= 8'h23;
            13'h0E3B: rddata <= 8'h23;
            13'h0E3C: rddata <= 8'hE5;
            13'h0E3D: rddata <= 8'hCD;
            13'h0E3E: rddata <= 8'hB3;
            13'h0E3F: rddata <= 8'h0E;
            13'h0E40: rddata <= 8'hE1;
            13'h0E41: rddata <= 8'h4E;
            13'h0E42: rddata <= 8'h23;
            13'h0E43: rddata <= 8'h46;
            13'h0E44: rddata <= 8'hCD;
            13'h0E45: rddata <= 8'h53;
            13'h0E46: rddata <= 8'h0E;
            13'h0E47: rddata <= 8'hE5;
            13'h0E48: rddata <= 8'h6F;
            13'h0E49: rddata <= 8'hCD;
            13'h0E4A: rddata <= 8'hBD;
            13'h0E4B: rddata <= 8'h0F;
            13'h0E4C: rddata <= 8'hD1;
            13'h0E4D: rddata <= 8'hC9;
            13'h0E4E: rddata <= 8'h3E;
            13'h0E4F: rddata <= 8'h01;
            13'h0E50: rddata <= 8'hCD;
            13'h0E51: rddata <= 8'hB3;
            13'h0E52: rddata <= 8'h0E;
            13'h0E53: rddata <= 8'h21;
            13'h0E54: rddata <= 8'hBD;
            13'h0E55: rddata <= 8'h38;
            13'h0E56: rddata <= 8'hE5;
            13'h0E57: rddata <= 8'h77;
            13'h0E58: rddata <= 8'h23;
            13'h0E59: rddata <= 8'h23;
            13'h0E5A: rddata <= 8'h73;
            13'h0E5B: rddata <= 8'h23;
            13'h0E5C: rddata <= 8'h72;
            13'h0E5D: rddata <= 8'hE1;
            13'h0E5E: rddata <= 8'hC9;
            13'h0E5F: rddata <= 8'h2B;
            13'h0E60: rddata <= 8'h06;
            13'h0E61: rddata <= 8'h22;
            13'h0E62: rddata <= 8'h50;
            13'h0E63: rddata <= 8'hE5;
            13'h0E64: rddata <= 8'h0E;
            13'h0E65: rddata <= 8'hFF;
            13'h0E66: rddata <= 8'h23;
            13'h0E67: rddata <= 8'h7E;
            13'h0E68: rddata <= 8'h0C;
            13'h0E69: rddata <= 8'hB7;
            13'h0E6A: rddata <= 8'h28;
            13'h0E6B: rddata <= 8'h06;
            13'h0E6C: rddata <= 8'hBA;
            13'h0E6D: rddata <= 8'h28;
            13'h0E6E: rddata <= 8'h03;
            13'h0E6F: rddata <= 8'hB8;
            13'h0E70: rddata <= 8'h20;
            13'h0E71: rddata <= 8'hF4;
            13'h0E72: rddata <= 8'hFE;
            13'h0E73: rddata <= 8'h22;
            13'h0E74: rddata <= 8'hCC;
            13'h0E75: rddata <= 8'h6B;
            13'h0E76: rddata <= 8'h06;
            13'h0E77: rddata <= 8'hE3;
            13'h0E78: rddata <= 8'h23;
            13'h0E79: rddata <= 8'hEB;
            13'h0E7A: rddata <= 8'h79;
            13'h0E7B: rddata <= 8'hCD;
            13'h0E7C: rddata <= 8'h53;
            13'h0E7D: rddata <= 8'h0E;
            13'h0E7E: rddata <= 8'h11;
            13'h0E7F: rddata <= 8'hBD;
            13'h0E80: rddata <= 8'h38;
            13'h0E81: rddata <= 8'h2A;
            13'h0E82: rddata <= 8'hAF;
            13'h0E83: rddata <= 8'h38;
            13'h0E84: rddata <= 8'h22;
            13'h0E85: rddata <= 8'hE4;
            13'h0E86: rddata <= 8'h38;
            13'h0E87: rddata <= 8'h3E;
            13'h0E88: rddata <= 8'h01;
            13'h0E89: rddata <= 8'h32;
            13'h0E8A: rddata <= 8'hAB;
            13'h0E8B: rddata <= 8'h38;
            13'h0E8C: rddata <= 8'hCD;
            13'h0E8D: rddata <= 8'h3D;
            13'h0E8E: rddata <= 8'h15;
            13'h0E8F: rddata <= 8'hE7;
            13'h0E90: rddata <= 8'h22;
            13'h0E91: rddata <= 8'hAF;
            13'h0E92: rddata <= 8'h38;
            13'h0E93: rddata <= 8'hE1;
            13'h0E94: rddata <= 8'h7E;
            13'h0E95: rddata <= 8'hC0;
            13'h0E96: rddata <= 8'h11;
            13'h0E97: rddata <= 8'h1E;
            13'h0E98: rddata <= 8'h00;
            13'h0E99: rddata <= 8'hC3;
            13'h0E9A: rddata <= 8'hDB;
            13'h0E9B: rddata <= 8'h03;
            13'h0E9C: rddata <= 8'h23;
            13'h0E9D: rddata <= 8'hCD;
            13'h0E9E: rddata <= 8'h5F;
            13'h0E9F: rddata <= 8'h0E;
            13'h0EA0: rddata <= 8'hCD;
            13'h0EA1: rddata <= 8'hC9;
            13'h0EA2: rddata <= 8'h0F;
            13'h0EA3: rddata <= 8'hCD;
            13'h0EA4: rddata <= 8'h31;
            13'h0EA5: rddata <= 8'h15;
            13'h0EA6: rddata <= 8'h1C;
            13'h0EA7: rddata <= 8'h1D;
            13'h0EA8: rddata <= 8'hC8;
            13'h0EA9: rddata <= 8'h0A;
            13'h0EAA: rddata <= 8'hDF;
            13'h0EAB: rddata <= 8'hFE;
            13'h0EAC: rddata <= 8'h0D;
            13'h0EAD: rddata <= 8'hCC;
            13'h0EAE: rddata <= 8'hF0;
            13'h0EAF: rddata <= 8'h19;
            13'h0EB0: rddata <= 8'h03;
            13'h0EB1: rddata <= 8'h18;
            13'h0EB2: rddata <= 8'hF4;
            13'h0EB3: rddata <= 8'hB7;
            13'h0EB4: rddata <= 8'h0E;
            13'h0EB5: rddata <= 8'hF1;
            13'h0EB6: rddata <= 8'hF5;
            13'h0EB7: rddata <= 8'h2A;
            13'h0EB8: rddata <= 8'h4B;
            13'h0EB9: rddata <= 8'h38;
            13'h0EBA: rddata <= 8'hEB;
            13'h0EBB: rddata <= 8'h2A;
            13'h0EBC: rddata <= 8'hC1;
            13'h0EBD: rddata <= 8'h38;
            13'h0EBE: rddata <= 8'h2F;
            13'h0EBF: rddata <= 8'h4F;
            13'h0EC0: rddata <= 8'h06;
            13'h0EC1: rddata <= 8'hFF;
            13'h0EC2: rddata <= 8'h09;
            13'h0EC3: rddata <= 8'h23;
            13'h0EC4: rddata <= 8'hE7;
            13'h0EC5: rddata <= 8'h38;
            13'h0EC6: rddata <= 8'h07;
            13'h0EC7: rddata <= 8'h22;
            13'h0EC8: rddata <= 8'hC1;
            13'h0EC9: rddata <= 8'h38;
            13'h0ECA: rddata <= 8'h23;
            13'h0ECB: rddata <= 8'hEB;
            13'h0ECC: rddata <= 8'hF1;
            13'h0ECD: rddata <= 8'hC9;
            13'h0ECE: rddata <= 8'hF1;
            13'h0ECF: rddata <= 8'h11;
            13'h0ED0: rddata <= 8'h1A;
            13'h0ED1: rddata <= 8'h00;
            13'h0ED2: rddata <= 8'hCA;
            13'h0ED3: rddata <= 8'hDB;
            13'h0ED4: rddata <= 8'h03;
            13'h0ED5: rddata <= 8'hBF;
            13'h0ED6: rddata <= 8'hF5;
            13'h0ED7: rddata <= 8'h01;
            13'h0ED8: rddata <= 8'hB5;
            13'h0ED9: rddata <= 8'h0E;
            13'h0EDA: rddata <= 8'hC5;
            13'h0EDB: rddata <= 8'h2A;
            13'h0EDC: rddata <= 8'hAD;
            13'h0EDD: rddata <= 8'h38;
            13'h0EDE: rddata <= 8'h22;
            13'h0EDF: rddata <= 8'hC1;
            13'h0EE0: rddata <= 8'h38;
            13'h0EE1: rddata <= 8'h21;
            13'h0EE2: rddata <= 8'h00;
            13'h0EE3: rddata <= 8'h00;
            13'h0EE4: rddata <= 8'hE5;
            13'h0EE5: rddata <= 8'h2A;
            13'h0EE6: rddata <= 8'hDA;
            13'h0EE7: rddata <= 8'h38;
            13'h0EE8: rddata <= 8'hE5;
            13'h0EE9: rddata <= 8'h21;
            13'h0EEA: rddata <= 8'hB1;
            13'h0EEB: rddata <= 8'h38;
            13'h0EEC: rddata <= 8'hED;
            13'h0EED: rddata <= 8'h5B;
            13'h0EEE: rddata <= 8'hAF;
            13'h0EEF: rddata <= 8'h38;
            13'h0EF0: rddata <= 8'hE7;
            13'h0EF1: rddata <= 8'h01;
            13'h0EF2: rddata <= 8'hEC;
            13'h0EF3: rddata <= 8'h0E;
            13'h0EF4: rddata <= 8'hC2;
            13'h0EF5: rddata <= 8'h32;
            13'h0EF6: rddata <= 8'h0F;
            13'h0EF7: rddata <= 8'h2A;
            13'h0EF8: rddata <= 8'hD6;
            13'h0EF9: rddata <= 8'h38;
            13'h0EFA: rddata <= 8'hED;
            13'h0EFB: rddata <= 8'h5B;
            13'h0EFC: rddata <= 8'hD8;
            13'h0EFD: rddata <= 8'h38;
            13'h0EFE: rddata <= 8'hE7;
            13'h0EFF: rddata <= 8'h28;
            13'h0F00: rddata <= 8'h0A;
            13'h0F01: rddata <= 8'h23;
            13'h0F02: rddata <= 8'h7E;
            13'h0F03: rddata <= 8'h23;
            13'h0F04: rddata <= 8'hB7;
            13'h0F05: rddata <= 8'hCD;
            13'h0F06: rddata <= 8'h35;
            13'h0F07: rddata <= 8'h0F;
            13'h0F08: rddata <= 8'h18;
            13'h0F09: rddata <= 8'hF0;
            13'h0F0A: rddata <= 8'hC1;
            13'h0F0B: rddata <= 8'hED;
            13'h0F0C: rddata <= 8'h5B;
            13'h0F0D: rddata <= 8'hDA;
            13'h0F0E: rddata <= 8'h38;
            13'h0F0F: rddata <= 8'hE7;
            13'h0F10: rddata <= 8'hCA;
            13'h0F11: rddata <= 8'h57;
            13'h0F12: rddata <= 8'h0F;
            13'h0F13: rddata <= 8'hCD;
            13'h0F14: rddata <= 8'h31;
            13'h0F15: rddata <= 8'h15;
            13'h0F16: rddata <= 8'h7A;
            13'h0F17: rddata <= 8'hE5;
            13'h0F18: rddata <= 8'h09;
            13'h0F19: rddata <= 8'hB7;
            13'h0F1A: rddata <= 8'hF2;
            13'h0F1B: rddata <= 8'h0A;
            13'h0F1C: rddata <= 8'h0F;
            13'h0F1D: rddata <= 8'h22;
            13'h0F1E: rddata <= 8'hC5;
            13'h0F1F: rddata <= 8'h38;
            13'h0F20: rddata <= 8'hE1;
            13'h0F21: rddata <= 8'h4E;
            13'h0F22: rddata <= 8'h06;
            13'h0F23: rddata <= 8'h00;
            13'h0F24: rddata <= 8'h09;
            13'h0F25: rddata <= 8'h09;
            13'h0F26: rddata <= 8'h23;
            13'h0F27: rddata <= 8'hEB;
            13'h0F28: rddata <= 8'h2A;
            13'h0F29: rddata <= 8'hC5;
            13'h0F2A: rddata <= 8'h38;
            13'h0F2B: rddata <= 8'hEB;
            13'h0F2C: rddata <= 8'hE7;
            13'h0F2D: rddata <= 8'h28;
            13'h0F2E: rddata <= 8'hDC;
            13'h0F2F: rddata <= 8'h01;
            13'h0F30: rddata <= 8'h27;
            13'h0F31: rddata <= 8'h0F;
            13'h0F32: rddata <= 8'hC5;
            13'h0F33: rddata <= 8'hF6;
            13'h0F34: rddata <= 8'h80;
            13'h0F35: rddata <= 8'h7E;
            13'h0F36: rddata <= 8'h23;
            13'h0F37: rddata <= 8'h23;
            13'h0F38: rddata <= 8'h5E;
            13'h0F39: rddata <= 8'h23;
            13'h0F3A: rddata <= 8'h56;
            13'h0F3B: rddata <= 8'h23;
            13'h0F3C: rddata <= 8'hF0;
            13'h0F3D: rddata <= 8'hB7;
            13'h0F3E: rddata <= 8'hC8;
            13'h0F3F: rddata <= 8'h44;
            13'h0F40: rddata <= 8'h4D;
            13'h0F41: rddata <= 8'h2A;
            13'h0F42: rddata <= 8'hC1;
            13'h0F43: rddata <= 8'h38;
            13'h0F44: rddata <= 8'hE7;
            13'h0F45: rddata <= 8'h60;
            13'h0F46: rddata <= 8'h69;
            13'h0F47: rddata <= 8'hD8;
            13'h0F48: rddata <= 8'hE1;
            13'h0F49: rddata <= 8'hE3;
            13'h0F4A: rddata <= 8'hE7;
            13'h0F4B: rddata <= 8'hE3;
            13'h0F4C: rddata <= 8'hE5;
            13'h0F4D: rddata <= 8'h60;
            13'h0F4E: rddata <= 8'h69;
            13'h0F4F: rddata <= 8'hD0;
            13'h0F50: rddata <= 8'hC1;
            13'h0F51: rddata <= 8'hF1;
            13'h0F52: rddata <= 8'hF1;
            13'h0F53: rddata <= 8'hE5;
            13'h0F54: rddata <= 8'hD5;
            13'h0F55: rddata <= 8'hC5;
            13'h0F56: rddata <= 8'hC9;
            13'h0F57: rddata <= 8'hD1;
            13'h0F58: rddata <= 8'hE1;
            13'h0F59: rddata <= 8'h7C;
            13'h0F5A: rddata <= 8'hB5;
            13'h0F5B: rddata <= 8'hC8;
            13'h0F5C: rddata <= 8'h2B;
            13'h0F5D: rddata <= 8'h46;
            13'h0F5E: rddata <= 8'h2B;
            13'h0F5F: rddata <= 8'h4E;
            13'h0F60: rddata <= 8'hE5;
            13'h0F61: rddata <= 8'h2B;
            13'h0F62: rddata <= 8'h2B;
            13'h0F63: rddata <= 8'h6E;
            13'h0F64: rddata <= 8'h26;
            13'h0F65: rddata <= 8'h00;
            13'h0F66: rddata <= 8'h09;
            13'h0F67: rddata <= 8'h50;
            13'h0F68: rddata <= 8'h59;
            13'h0F69: rddata <= 8'h2B;
            13'h0F6A: rddata <= 8'h44;
            13'h0F6B: rddata <= 8'h4D;
            13'h0F6C: rddata <= 8'h2A;
            13'h0F6D: rddata <= 8'hC1;
            13'h0F6E: rddata <= 8'h38;
            13'h0F6F: rddata <= 8'hCD;
            13'h0F70: rddata <= 8'h95;
            13'h0F71: rddata <= 8'h0B;
            13'h0F72: rddata <= 8'hE1;
            13'h0F73: rddata <= 8'h71;
            13'h0F74: rddata <= 8'h23;
            13'h0F75: rddata <= 8'h70;
            13'h0F76: rddata <= 8'h60;
            13'h0F77: rddata <= 8'h69;
            13'h0F78: rddata <= 8'h2B;
            13'h0F79: rddata <= 8'hC3;
            13'h0F7A: rddata <= 8'hDE;
            13'h0F7B: rddata <= 8'h0E;
            13'h0F7C: rddata <= 8'hC5;
            13'h0F7D: rddata <= 8'hE5;
            13'h0F7E: rddata <= 8'h2A;
            13'h0F7F: rddata <= 8'hE4;
            13'h0F80: rddata <= 8'h38;
            13'h0F81: rddata <= 8'hE3;
            13'h0F82: rddata <= 8'hCD;
            13'h0F83: rddata <= 8'hFD;
            13'h0F84: rddata <= 8'h09;
            13'h0F85: rddata <= 8'hE3;
            13'h0F86: rddata <= 8'hCD;
            13'h0F87: rddata <= 8'h76;
            13'h0F88: rddata <= 8'h09;
            13'h0F89: rddata <= 8'h7E;
            13'h0F8A: rddata <= 8'hE5;
            13'h0F8B: rddata <= 8'h2A;
            13'h0F8C: rddata <= 8'hE4;
            13'h0F8D: rddata <= 8'h38;
            13'h0F8E: rddata <= 8'hE5;
            13'h0F8F: rddata <= 8'h86;
            13'h0F90: rddata <= 8'h11;
            13'h0F91: rddata <= 8'h1C;
            13'h0F92: rddata <= 8'h00;
            13'h0F93: rddata <= 8'hDA;
            13'h0F94: rddata <= 8'hDB;
            13'h0F95: rddata <= 8'h03;
            13'h0F96: rddata <= 8'hCD;
            13'h0F97: rddata <= 8'h50;
            13'h0F98: rddata <= 8'h0E;
            13'h0F99: rddata <= 8'hD1;
            13'h0F9A: rddata <= 8'hCD;
            13'h0F9B: rddata <= 8'hCD;
            13'h0F9C: rddata <= 8'h0F;
            13'h0F9D: rddata <= 8'hE3;
            13'h0F9E: rddata <= 8'hCD;
            13'h0F9F: rddata <= 8'hCC;
            13'h0FA0: rddata <= 8'h0F;
            13'h0FA1: rddata <= 8'hE5;
            13'h0FA2: rddata <= 8'h2A;
            13'h0FA3: rddata <= 8'hBF;
            13'h0FA4: rddata <= 8'h38;
            13'h0FA5: rddata <= 8'hEB;
            13'h0FA6: rddata <= 8'hCD;
            13'h0FA7: rddata <= 8'hB4;
            13'h0FA8: rddata <= 8'h0F;
            13'h0FA9: rddata <= 8'hCD;
            13'h0FAA: rddata <= 8'hB4;
            13'h0FAB: rddata <= 8'h0F;
            13'h0FAC: rddata <= 8'h21;
            13'h0FAD: rddata <= 8'h91;
            13'h0FAE: rddata <= 8'h09;
            13'h0FAF: rddata <= 8'hE3;
            13'h0FB0: rddata <= 8'hE5;
            13'h0FB1: rddata <= 8'hC3;
            13'h0FB2: rddata <= 8'h7E;
            13'h0FB3: rddata <= 8'h0E;
            13'h0FB4: rddata <= 8'hE1;
            13'h0FB5: rddata <= 8'hE3;
            13'h0FB6: rddata <= 8'h7E;
            13'h0FB7: rddata <= 8'h23;
            13'h0FB8: rddata <= 8'h23;
            13'h0FB9: rddata <= 8'h4E;
            13'h0FBA: rddata <= 8'h23;
            13'h0FBB: rddata <= 8'h46;
            13'h0FBC: rddata <= 8'h6F;
            13'h0FBD: rddata <= 8'h2C;
            13'h0FBE: rddata <= 8'h2D;
            13'h0FBF: rddata <= 8'hC8;
            13'h0FC0: rddata <= 8'h0A;
            13'h0FC1: rddata <= 8'h12;
            13'h0FC2: rddata <= 8'h03;
            13'h0FC3: rddata <= 8'h13;
            13'h0FC4: rddata <= 8'h18;
            13'h0FC5: rddata <= 8'hF8;
            13'h0FC6: rddata <= 8'hCD;
            13'h0FC7: rddata <= 8'h76;
            13'h0FC8: rddata <= 8'h09;
            13'h0FC9: rddata <= 8'h2A;
            13'h0FCA: rddata <= 8'hE4;
            13'h0FCB: rddata <= 8'h38;
            13'h0FCC: rddata <= 8'hEB;
            13'h0FCD: rddata <= 8'hCD;
            13'h0FCE: rddata <= 8'hE4;
            13'h0FCF: rddata <= 8'h0F;
            13'h0FD0: rddata <= 8'hEB;
            13'h0FD1: rddata <= 8'hC0;
            13'h0FD2: rddata <= 8'hD5;
            13'h0FD3: rddata <= 8'h50;
            13'h0FD4: rddata <= 8'h59;
            13'h0FD5: rddata <= 8'h1B;
            13'h0FD6: rddata <= 8'h4E;
            13'h0FD7: rddata <= 8'h2A;
            13'h0FD8: rddata <= 8'hC1;
            13'h0FD9: rddata <= 8'h38;
            13'h0FDA: rddata <= 8'hE7;
            13'h0FDB: rddata <= 8'h20;
            13'h0FDC: rddata <= 8'h05;
            13'h0FDD: rddata <= 8'h47;
            13'h0FDE: rddata <= 8'h09;
            13'h0FDF: rddata <= 8'h22;
            13'h0FE0: rddata <= 8'hC1;
            13'h0FE1: rddata <= 8'h38;
            13'h0FE2: rddata <= 8'hE1;
            13'h0FE3: rddata <= 8'hC9;
            13'h0FE4: rddata <= 8'h2A;
            13'h0FE5: rddata <= 8'hAF;
            13'h0FE6: rddata <= 8'h38;
            13'h0FE7: rddata <= 8'h2B;
            13'h0FE8: rddata <= 8'h46;
            13'h0FE9: rddata <= 8'h2B;
            13'h0FEA: rddata <= 8'h4E;
            13'h0FEB: rddata <= 8'h2B;
            13'h0FEC: rddata <= 8'h2B;
            13'h0FED: rddata <= 8'hE7;
            13'h0FEE: rddata <= 8'hC0;
            13'h0FEF: rddata <= 8'h22;
            13'h0FF0: rddata <= 8'hAF;
            13'h0FF1: rddata <= 8'h38;
            13'h0FF2: rddata <= 8'hC9;
            13'h0FF3: rddata <= 8'h01;
            13'h0FF4: rddata <= 8'h36;
            13'h0FF5: rddata <= 8'h0B;
            13'h0FF6: rddata <= 8'hC5;
            13'h0FF7: rddata <= 8'hCD;
            13'h0FF8: rddata <= 8'hC6;
            13'h0FF9: rddata <= 8'h0F;
            13'h0FFA: rddata <= 8'hAF;
            13'h0FFB: rddata <= 8'h57;
            13'h0FFC: rddata <= 8'h32;
            13'h0FFD: rddata <= 8'hAB;
            13'h0FFE: rddata <= 8'h38;
            13'h0FFF: rddata <= 8'h7E;
            13'h1000: rddata <= 8'hB7;
            13'h1001: rddata <= 8'hC9;
            13'h1002: rddata <= 8'h01;
            13'h1003: rddata <= 8'h36;
            13'h1004: rddata <= 8'h0B;
            13'h1005: rddata <= 8'hC5;
            13'h1006: rddata <= 8'hCD;
            13'h1007: rddata <= 8'hF7;
            13'h1008: rddata <= 8'h0F;
            13'h1009: rddata <= 8'hCA;
            13'h100A: rddata <= 8'h97;
            13'h100B: rddata <= 8'h06;
            13'h100C: rddata <= 8'h23;
            13'h100D: rddata <= 8'h23;
            13'h100E: rddata <= 8'h5E;
            13'h100F: rddata <= 8'h23;
            13'h1010: rddata <= 8'h56;
            13'h1011: rddata <= 8'h1A;
            13'h1012: rddata <= 8'hC9;
            13'h1013: rddata <= 8'hCD;
            13'h1014: rddata <= 8'h4E;
            13'h1015: rddata <= 8'h0E;
            13'h1016: rddata <= 8'hCD;
            13'h1017: rddata <= 8'h57;
            13'h1018: rddata <= 8'h0B;
            13'h1019: rddata <= 8'h2A;
            13'h101A: rddata <= 8'hBF;
            13'h101B: rddata <= 8'h38;
            13'h101C: rddata <= 8'h73;
            13'h101D: rddata <= 8'hC1;
            13'h101E: rddata <= 8'hC3;
            13'h101F: rddata <= 8'h7E;
            13'h1020: rddata <= 8'h0E;
            13'h1021: rddata <= 8'hCD;
            13'h1022: rddata <= 8'hA0;
            13'h1023: rddata <= 8'h10;
            13'h1024: rddata <= 8'hAF;
            13'h1025: rddata <= 8'hE3;
            13'h1026: rddata <= 8'h4F;
            13'h1027: rddata <= 8'hE5;
            13'h1028: rddata <= 8'h7E;
            13'h1029: rddata <= 8'hB8;
            13'h102A: rddata <= 8'h38;
            13'h102B: rddata <= 8'h02;
            13'h102C: rddata <= 8'h78;
            13'h102D: rddata <= 8'h11;
            13'h102E: rddata <= 8'h0E;
            13'h102F: rddata <= 8'h00;
            13'h1030: rddata <= 8'hC5;
            13'h1031: rddata <= 8'hCD;
            13'h1032: rddata <= 8'hB3;
            13'h1033: rddata <= 8'h0E;
            13'h1034: rddata <= 8'hC1;
            13'h1035: rddata <= 8'hE1;
            13'h1036: rddata <= 8'hE5;
            13'h1037: rddata <= 8'h23;
            13'h1038: rddata <= 8'h23;
            13'h1039: rddata <= 8'h46;
            13'h103A: rddata <= 8'h23;
            13'h103B: rddata <= 8'h66;
            13'h103C: rddata <= 8'h68;
            13'h103D: rddata <= 8'h06;
            13'h103E: rddata <= 8'h00;
            13'h103F: rddata <= 8'h09;
            13'h1040: rddata <= 8'h44;
            13'h1041: rddata <= 8'h4D;
            13'h1042: rddata <= 8'hCD;
            13'h1043: rddata <= 8'h53;
            13'h1044: rddata <= 8'h0E;
            13'h1045: rddata <= 8'h6F;
            13'h1046: rddata <= 8'hCD;
            13'h1047: rddata <= 8'hBD;
            13'h1048: rddata <= 8'h0F;
            13'h1049: rddata <= 8'hD1;
            13'h104A: rddata <= 8'hCD;
            13'h104B: rddata <= 8'hCD;
            13'h104C: rddata <= 8'h0F;
            13'h104D: rddata <= 8'hC3;
            13'h104E: rddata <= 8'h7E;
            13'h104F: rddata <= 8'h0E;
            13'h1050: rddata <= 8'hCD;
            13'h1051: rddata <= 8'hA0;
            13'h1052: rddata <= 8'h10;
            13'h1053: rddata <= 8'hD1;
            13'h1054: rddata <= 8'hD5;
            13'h1055: rddata <= 8'h1A;
            13'h1056: rddata <= 8'h90;
            13'h1057: rddata <= 8'h18;
            13'h1058: rddata <= 8'hCC;
            13'h1059: rddata <= 8'hEB;
            13'h105A: rddata <= 8'h7E;
            13'h105B: rddata <= 8'hCD;
            13'h105C: rddata <= 8'hA3;
            13'h105D: rddata <= 8'h10;
            13'h105E: rddata <= 8'h04;
            13'h105F: rddata <= 8'h05;
            13'h1060: rddata <= 8'hCA;
            13'h1061: rddata <= 8'h97;
            13'h1062: rddata <= 8'h06;
            13'h1063: rddata <= 8'hC5;
            13'h1064: rddata <= 8'h1E;
            13'h1065: rddata <= 8'hFF;
            13'h1066: rddata <= 8'hFE;
            13'h1067: rddata <= 8'h29;
            13'h1068: rddata <= 8'h28;
            13'h1069: rddata <= 8'h05;
            13'h106A: rddata <= 8'hCF;
            13'h106B: rddata <= 8'h2C;
            13'h106C: rddata <= 8'hCD;
            13'h106D: rddata <= 8'h54;
            13'h106E: rddata <= 8'h0B;
            13'h106F: rddata <= 8'hCF;
            13'h1070: rddata <= 8'h29;
            13'h1071: rddata <= 8'hF1;
            13'h1072: rddata <= 8'hE3;
            13'h1073: rddata <= 8'h01;
            13'h1074: rddata <= 8'h27;
            13'h1075: rddata <= 8'h10;
            13'h1076: rddata <= 8'hC5;
            13'h1077: rddata <= 8'h3D;
            13'h1078: rddata <= 8'hBE;
            13'h1079: rddata <= 8'h06;
            13'h107A: rddata <= 8'h00;
            13'h107B: rddata <= 8'hD0;
            13'h107C: rddata <= 8'h4F;
            13'h107D: rddata <= 8'h7E;
            13'h107E: rddata <= 8'h91;
            13'h107F: rddata <= 8'hBB;
            13'h1080: rddata <= 8'h47;
            13'h1081: rddata <= 8'hD8;
            13'h1082: rddata <= 8'h43;
            13'h1083: rddata <= 8'hC9;
            13'h1084: rddata <= 8'hCD;
            13'h1085: rddata <= 8'hF7;
            13'h1086: rddata <= 8'h0F;
            13'h1087: rddata <= 8'hCA;
            13'h1088: rddata <= 8'hC3;
            13'h1089: rddata <= 8'h12;
            13'h108A: rddata <= 8'h5F;
            13'h108B: rddata <= 8'h23;
            13'h108C: rddata <= 8'h23;
            13'h108D: rddata <= 8'h7E;
            13'h108E: rddata <= 8'h23;
            13'h108F: rddata <= 8'h66;
            13'h1090: rddata <= 8'h6F;
            13'h1091: rddata <= 8'hE5;
            13'h1092: rddata <= 8'h19;
            13'h1093: rddata <= 8'h46;
            13'h1094: rddata <= 8'h72;
            13'h1095: rddata <= 8'hE3;
            13'h1096: rddata <= 8'hC5;
            13'h1097: rddata <= 8'h2B;
            13'h1098: rddata <= 8'hD7;
            13'h1099: rddata <= 8'hCD;
            13'h109A: rddata <= 8'hE5;
            13'h109B: rddata <= 8'h15;
            13'h109C: rddata <= 8'hC1;
            13'h109D: rddata <= 8'hE1;
            13'h109E: rddata <= 8'h70;
            13'h109F: rddata <= 8'hC9;
            13'h10A0: rddata <= 8'hEB;
            13'h10A1: rddata <= 8'hCF;
            13'h10A2: rddata <= 8'h29;
            13'h10A3: rddata <= 8'hC1;
            13'h10A4: rddata <= 8'hD1;
            13'h10A5: rddata <= 8'hC5;
            13'h10A6: rddata <= 8'h43;
            13'h10A7: rddata <= 8'hC9;
            13'h10A8: rddata <= 8'h2A;
            13'h10A9: rddata <= 8'hDA;
            13'h10AA: rddata <= 8'h38;
            13'h10AB: rddata <= 8'hEB;
            13'h10AC: rddata <= 8'h21;
            13'h10AD: rddata <= 8'h00;
            13'h10AE: rddata <= 8'h00;
            13'h10AF: rddata <= 8'h39;
            13'h10B0: rddata <= 8'h3A;
            13'h10B1: rddata <= 8'hAB;
            13'h10B2: rddata <= 8'h38;
            13'h10B3: rddata <= 8'hB7;
            13'h10B4: rddata <= 8'hCA;
            13'h10B5: rddata <= 8'h1C;
            13'h10B6: rddata <= 8'h0B;
            13'h10B7: rddata <= 8'hCD;
            13'h10B8: rddata <= 8'hC9;
            13'h10B9: rddata <= 8'h0F;
            13'h10BA: rddata <= 8'hCD;
            13'h10BB: rddata <= 8'hDB;
            13'h10BC: rddata <= 8'h0E;
            13'h10BD: rddata <= 8'hED;
            13'h10BE: rddata <= 8'h5B;
            13'h10BF: rddata <= 8'h4B;
            13'h10C0: rddata <= 8'h38;
            13'h10C1: rddata <= 8'h2A;
            13'h10C2: rddata <= 8'hC1;
            13'h10C3: rddata <= 8'h38;
            13'h10C4: rddata <= 8'hC3;
            13'h10C5: rddata <= 8'h1C;
            13'h10C6: rddata <= 8'h0B;
            13'h10C7: rddata <= 8'h2B;
            13'h10C8: rddata <= 8'hD7;
            13'h10C9: rddata <= 8'hC8;
            13'h10CA: rddata <= 8'hCF;
            13'h10CB: rddata <= 8'h2C;
            13'h10CC: rddata <= 8'h01;
            13'h10CD: rddata <= 8'hC7;
            13'h10CE: rddata <= 8'h10;
            13'h10CF: rddata <= 8'hC5;
            13'h10D0: rddata <= 8'hF6;
            13'h10D1: rddata <= 8'hAF;
            13'h10D2: rddata <= 8'h32;
            13'h10D3: rddata <= 8'hAA;
            13'h10D4: rddata <= 8'h38;
            13'h10D5: rddata <= 8'h4E;
            13'h10D6: rddata <= 8'hCD;
            13'h10D7: rddata <= 8'hC5;
            13'h10D8: rddata <= 8'h0C;
            13'h10D9: rddata <= 8'hDA;
            13'h10DA: rddata <= 8'hC4;
            13'h10DB: rddata <= 8'h03;
            13'h10DC: rddata <= 8'hAF;
            13'h10DD: rddata <= 8'h47;
            13'h10DE: rddata <= 8'h32;
            13'h10DF: rddata <= 8'hAB;
            13'h10E0: rddata <= 8'h38;
            13'h10E1: rddata <= 8'hD7;
            13'h10E2: rddata <= 8'h38;
            13'h10E3: rddata <= 8'h05;
            13'h10E4: rddata <= 8'hCD;
            13'h10E5: rddata <= 8'hC6;
            13'h10E6: rddata <= 8'h0C;
            13'h10E7: rddata <= 8'h38;
            13'h10E8: rddata <= 8'h09;
            13'h10E9: rddata <= 8'h47;
            13'h10EA: rddata <= 8'hD7;
            13'h10EB: rddata <= 8'h38;
            13'h10EC: rddata <= 8'hFD;
            13'h10ED: rddata <= 8'hCD;
            13'h10EE: rddata <= 8'hC6;
            13'h10EF: rddata <= 8'h0C;
            13'h10F0: rddata <= 8'h30;
            13'h10F1: rddata <= 8'hF8;
            13'h10F2: rddata <= 8'hD6;
            13'h10F3: rddata <= 8'h24;
            13'h10F4: rddata <= 8'h20;
            13'h10F5: rddata <= 8'h08;
            13'h10F6: rddata <= 8'h3C;
            13'h10F7: rddata <= 8'h32;
            13'h10F8: rddata <= 8'hAB;
            13'h10F9: rddata <= 8'h38;
            13'h10FA: rddata <= 8'h0F;
            13'h10FB: rddata <= 8'h80;
            13'h10FC: rddata <= 8'h47;
            13'h10FD: rddata <= 8'hD7;
            13'h10FE: rddata <= 8'h3A;
            13'h10FF: rddata <= 8'hCB;
            13'h1100: rddata <= 8'h38;
            13'h1101: rddata <= 8'h3D;
            13'h1102: rddata <= 8'hCA;
            13'h1103: rddata <= 8'hA0;
            13'h1104: rddata <= 8'h11;
            13'h1105: rddata <= 8'hF2;
            13'h1106: rddata <= 8'h0E;
            13'h1107: rddata <= 8'h11;
            13'h1108: rddata <= 8'h7E;
            13'h1109: rddata <= 8'hD6;
            13'h110A: rddata <= 8'h28;
            13'h110B: rddata <= 8'hCA;
            13'h110C: rddata <= 8'h7A;
            13'h110D: rddata <= 8'h11;
            13'h110E: rddata <= 8'hAF;
            13'h110F: rddata <= 8'h32;
            13'h1110: rddata <= 8'hCB;
            13'h1111: rddata <= 8'h38;
            13'h1112: rddata <= 8'hE5;
            13'h1113: rddata <= 8'h50;
            13'h1114: rddata <= 8'h59;
            13'h1115: rddata <= 8'h2A;
            13'h1116: rddata <= 8'hDE;
            13'h1117: rddata <= 8'h38;
            13'h1118: rddata <= 8'hE7;
            13'h1119: rddata <= 8'h11;
            13'h111A: rddata <= 8'hE0;
            13'h111B: rddata <= 8'h38;
            13'h111C: rddata <= 8'hCA;
            13'h111D: rddata <= 8'h1A;
            13'h111E: rddata <= 8'h14;
            13'h111F: rddata <= 8'h2A;
            13'h1120: rddata <= 8'hD8;
            13'h1121: rddata <= 8'h38;
            13'h1122: rddata <= 8'hEB;
            13'h1123: rddata <= 8'h2A;
            13'h1124: rddata <= 8'hD6;
            13'h1125: rddata <= 8'h38;
            13'h1126: rddata <= 8'hE7;
            13'h1127: rddata <= 8'hCA;
            13'h1128: rddata <= 8'h3D;
            13'h1129: rddata <= 8'h11;
            13'h112A: rddata <= 8'h79;
            13'h112B: rddata <= 8'h96;
            13'h112C: rddata <= 8'h23;
            13'h112D: rddata <= 8'hC2;
            13'h112E: rddata <= 8'h32;
            13'h112F: rddata <= 8'h11;
            13'h1130: rddata <= 8'h78;
            13'h1131: rddata <= 8'h96;
            13'h1132: rddata <= 8'h23;
            13'h1133: rddata <= 8'hCA;
            13'h1134: rddata <= 8'h6C;
            13'h1135: rddata <= 8'h11;
            13'h1136: rddata <= 8'h23;
            13'h1137: rddata <= 8'h23;
            13'h1138: rddata <= 8'h23;
            13'h1139: rddata <= 8'h23;
            13'h113A: rddata <= 8'hC3;
            13'h113B: rddata <= 8'h26;
            13'h113C: rddata <= 8'h11;
            13'h113D: rddata <= 8'hE1;
            13'h113E: rddata <= 8'hE3;
            13'h113F: rddata <= 8'hD5;
            13'h1140: rddata <= 8'h11;
            13'h1141: rddata <= 8'h51;
            13'h1142: rddata <= 8'h0A;
            13'h1143: rddata <= 8'hE7;
            13'h1144: rddata <= 8'hD1;
            13'h1145: rddata <= 8'hCA;
            13'h1146: rddata <= 8'h6F;
            13'h1147: rddata <= 8'h11;
            13'h1148: rddata <= 8'hE3;
            13'h1149: rddata <= 8'hE5;
            13'h114A: rddata <= 8'hC5;
            13'h114B: rddata <= 8'h01;
            13'h114C: rddata <= 8'h06;
            13'h114D: rddata <= 8'h00;
            13'h114E: rddata <= 8'h2A;
            13'h114F: rddata <= 8'hDA;
            13'h1150: rddata <= 8'h38;
            13'h1151: rddata <= 8'hE5;
            13'h1152: rddata <= 8'h09;
            13'h1153: rddata <= 8'hC1;
            13'h1154: rddata <= 8'hE5;
            13'h1155: rddata <= 8'hCD;
            13'h1156: rddata <= 8'h92;
            13'h1157: rddata <= 8'h0B;
            13'h1158: rddata <= 8'hE1;
            13'h1159: rddata <= 8'h22;
            13'h115A: rddata <= 8'hDA;
            13'h115B: rddata <= 8'h38;
            13'h115C: rddata <= 8'h60;
            13'h115D: rddata <= 8'h69;
            13'h115E: rddata <= 8'h22;
            13'h115F: rddata <= 8'hD8;
            13'h1160: rddata <= 8'h38;
            13'h1161: rddata <= 8'h2B;
            13'h1162: rddata <= 8'h36;
            13'h1163: rddata <= 8'h00;
            13'h1164: rddata <= 8'hE7;
            13'h1165: rddata <= 8'h20;
            13'h1166: rddata <= 8'hFA;
            13'h1167: rddata <= 8'hD1;
            13'h1168: rddata <= 8'h73;
            13'h1169: rddata <= 8'h23;
            13'h116A: rddata <= 8'h72;
            13'h116B: rddata <= 8'h23;
            13'h116C: rddata <= 8'hEB;
            13'h116D: rddata <= 8'hE1;
            13'h116E: rddata <= 8'hC9;
            13'h116F: rddata <= 8'h32;
            13'h1170: rddata <= 8'hE7;
            13'h1171: rddata <= 8'h38;
            13'h1172: rddata <= 8'h21;
            13'h1173: rddata <= 8'h6D;
            13'h1174: rddata <= 8'h03;
            13'h1175: rddata <= 8'h22;
            13'h1176: rddata <= 8'hE4;
            13'h1177: rddata <= 8'h38;
            13'h1178: rddata <= 8'hE1;
            13'h1179: rddata <= 8'hC9;
            13'h117A: rddata <= 8'hE5;
            13'h117B: rddata <= 8'h2A;
            13'h117C: rddata <= 8'hAA;
            13'h117D: rddata <= 8'h38;
            13'h117E: rddata <= 8'hE3;
            13'h117F: rddata <= 8'h57;
            13'h1180: rddata <= 8'hD5;
            13'h1181: rddata <= 8'hC5;
            13'h1182: rddata <= 8'hCD;
            13'h1183: rddata <= 8'h7A;
            13'h1184: rddata <= 8'h06;
            13'h1185: rddata <= 8'hC1;
            13'h1186: rddata <= 8'hF1;
            13'h1187: rddata <= 8'hEB;
            13'h1188: rddata <= 8'hE3;
            13'h1189: rddata <= 8'hE5;
            13'h118A: rddata <= 8'hEB;
            13'h118B: rddata <= 8'h3C;
            13'h118C: rddata <= 8'h57;
            13'h118D: rddata <= 8'h7E;
            13'h118E: rddata <= 8'hFE;
            13'h118F: rddata <= 8'h2C;
            13'h1190: rddata <= 8'hCA;
            13'h1191: rddata <= 8'h80;
            13'h1192: rddata <= 8'h11;
            13'h1193: rddata <= 8'hCF;
            13'h1194: rddata <= 8'h29;
            13'h1195: rddata <= 8'h22;
            13'h1196: rddata <= 8'hD0;
            13'h1197: rddata <= 8'h38;
            13'h1198: rddata <= 8'hE1;
            13'h1199: rddata <= 8'h22;
            13'h119A: rddata <= 8'hAA;
            13'h119B: rddata <= 8'h38;
            13'h119C: rddata <= 8'h1E;
            13'h119D: rddata <= 8'h00;
            13'h119E: rddata <= 8'hD5;
            13'h119F: rddata <= 8'h11;
            13'h11A0: rddata <= 8'hE5;
            13'h11A1: rddata <= 8'hF5;
            13'h11A2: rddata <= 8'h2A;
            13'h11A3: rddata <= 8'hD8;
            13'h11A4: rddata <= 8'h38;
            13'h11A5: rddata <= 8'h3E;
            13'h11A6: rddata <= 8'h19;
            13'h11A7: rddata <= 8'hED;
            13'h11A8: rddata <= 8'h5B;
            13'h11A9: rddata <= 8'hDA;
            13'h11AA: rddata <= 8'h38;
            13'h11AB: rddata <= 8'hE7;
            13'h11AC: rddata <= 8'h28;
            13'h11AD: rddata <= 8'h25;
            13'h11AE: rddata <= 8'h7E;
            13'h11AF: rddata <= 8'h23;
            13'h11B0: rddata <= 8'hB9;
            13'h11B1: rddata <= 8'h20;
            13'h11B2: rddata <= 8'h02;
            13'h11B3: rddata <= 8'h7E;
            13'h11B4: rddata <= 8'hB8;
            13'h11B5: rddata <= 8'h23;
            13'h11B6: rddata <= 8'h5E;
            13'h11B7: rddata <= 8'h23;
            13'h11B8: rddata <= 8'h56;
            13'h11B9: rddata <= 8'h23;
            13'h11BA: rddata <= 8'h20;
            13'h11BB: rddata <= 8'hEA;
            13'h11BC: rddata <= 8'h3A;
            13'h11BD: rddata <= 8'hAA;
            13'h11BE: rddata <= 8'h38;
            13'h11BF: rddata <= 8'hB7;
            13'h11C0: rddata <= 8'hC2;
            13'h11C1: rddata <= 8'hCD;
            13'h11C2: rddata <= 8'h03;
            13'h11C3: rddata <= 8'hF1;
            13'h11C4: rddata <= 8'h44;
            13'h11C5: rddata <= 8'h4D;
            13'h11C6: rddata <= 8'hCA;
            13'h11C7: rddata <= 8'h1A;
            13'h11C8: rddata <= 8'h14;
            13'h11C9: rddata <= 8'h96;
            13'h11CA: rddata <= 8'hCA;
            13'h11CB: rddata <= 8'h2B;
            13'h11CC: rddata <= 8'h12;
            13'h11CD: rddata <= 8'h11;
            13'h11CE: rddata <= 8'h10;
            13'h11CF: rddata <= 8'h00;
            13'h11D0: rddata <= 8'hC3;
            13'h11D1: rddata <= 8'hDB;
            13'h11D2: rddata <= 8'h03;
            13'h11D3: rddata <= 8'h11;
            13'h11D4: rddata <= 8'h04;
            13'h11D5: rddata <= 8'h00;
            13'h11D6: rddata <= 8'hF1;
            13'h11D7: rddata <= 8'hCA;
            13'h11D8: rddata <= 8'h97;
            13'h11D9: rddata <= 8'h06;
            13'h11DA: rddata <= 8'h71;
            13'h11DB: rddata <= 8'h23;
            13'h11DC: rddata <= 8'h70;
            13'h11DD: rddata <= 8'h23;
            13'h11DE: rddata <= 8'h4F;
            13'h11DF: rddata <= 8'hCD;
            13'h11E0: rddata <= 8'hA0;
            13'h11E1: rddata <= 8'h0B;
            13'h11E2: rddata <= 8'h23;
            13'h11E3: rddata <= 8'h23;
            13'h11E4: rddata <= 8'h22;
            13'h11E5: rddata <= 8'hC3;
            13'h11E6: rddata <= 8'h38;
            13'h11E7: rddata <= 8'h71;
            13'h11E8: rddata <= 8'h23;
            13'h11E9: rddata <= 8'h3A;
            13'h11EA: rddata <= 8'hAA;
            13'h11EB: rddata <= 8'h38;
            13'h11EC: rddata <= 8'h17;
            13'h11ED: rddata <= 8'h79;
            13'h11EE: rddata <= 8'h01;
            13'h11EF: rddata <= 8'h0B;
            13'h11F0: rddata <= 8'h00;
            13'h11F1: rddata <= 8'h30;
            13'h11F2: rddata <= 8'h02;
            13'h11F3: rddata <= 8'hC1;
            13'h11F4: rddata <= 8'h03;
            13'h11F5: rddata <= 8'h71;
            13'h11F6: rddata <= 8'hF5;
            13'h11F7: rddata <= 8'h23;
            13'h11F8: rddata <= 8'h70;
            13'h11F9: rddata <= 8'h23;
            13'h11FA: rddata <= 8'hE5;
            13'h11FB: rddata <= 8'hCD;
            13'h11FC: rddata <= 8'hCA;
            13'h11FD: rddata <= 8'h15;
            13'h11FE: rddata <= 8'hEB;
            13'h11FF: rddata <= 8'hE1;
            13'h1200: rddata <= 8'hF1;
            13'h1201: rddata <= 8'h3D;
            13'h1202: rddata <= 8'h20;
            13'h1203: rddata <= 8'hEA;
            13'h1204: rddata <= 8'hF5;
            13'h1205: rddata <= 8'h42;
            13'h1206: rddata <= 8'h4B;
            13'h1207: rddata <= 8'hEB;
            13'h1208: rddata <= 8'h19;
            13'h1209: rddata <= 8'hDA;
            13'h120A: rddata <= 8'hB7;
            13'h120B: rddata <= 8'h0B;
            13'h120C: rddata <= 8'hCD;
            13'h120D: rddata <= 8'hA9;
            13'h120E: rddata <= 8'h0B;
            13'h120F: rddata <= 8'h22;
            13'h1210: rddata <= 8'hDA;
            13'h1211: rddata <= 8'h38;
            13'h1212: rddata <= 8'h2B;
            13'h1213: rddata <= 8'h36;
            13'h1214: rddata <= 8'h00;
            13'h1215: rddata <= 8'hE7;
            13'h1216: rddata <= 8'h20;
            13'h1217: rddata <= 8'hFA;
            13'h1218: rddata <= 8'h03;
            13'h1219: rddata <= 8'h57;
            13'h121A: rddata <= 8'h2A;
            13'h121B: rddata <= 8'hC3;
            13'h121C: rddata <= 8'h38;
            13'h121D: rddata <= 8'h5E;
            13'h121E: rddata <= 8'hEB;
            13'h121F: rddata <= 8'h29;
            13'h1220: rddata <= 8'h09;
            13'h1221: rddata <= 8'hEB;
            13'h1222: rddata <= 8'h2B;
            13'h1223: rddata <= 8'h2B;
            13'h1224: rddata <= 8'h73;
            13'h1225: rddata <= 8'h23;
            13'h1226: rddata <= 8'h72;
            13'h1227: rddata <= 8'h23;
            13'h1228: rddata <= 8'hF1;
            13'h1229: rddata <= 8'h38;
            13'h122A: rddata <= 8'h21;
            13'h122B: rddata <= 8'h47;
            13'h122C: rddata <= 8'h4F;
            13'h122D: rddata <= 8'h7E;
            13'h122E: rddata <= 8'h23;
            13'h122F: rddata <= 8'h16;
            13'h1230: rddata <= 8'hE1;
            13'h1231: rddata <= 8'h5E;
            13'h1232: rddata <= 8'h23;
            13'h1233: rddata <= 8'h56;
            13'h1234: rddata <= 8'h23;
            13'h1235: rddata <= 8'hE3;
            13'h1236: rddata <= 8'hF5;
            13'h1237: rddata <= 8'hE7;
            13'h1238: rddata <= 8'hD2;
            13'h1239: rddata <= 8'hCD;
            13'h123A: rddata <= 8'h11;
            13'h123B: rddata <= 8'hE5;
            13'h123C: rddata <= 8'hCD;
            13'h123D: rddata <= 8'hCA;
            13'h123E: rddata <= 8'h15;
            13'h123F: rddata <= 8'hD1;
            13'h1240: rddata <= 8'h19;
            13'h1241: rddata <= 8'hF1;
            13'h1242: rddata <= 8'h3D;
            13'h1243: rddata <= 8'h44;
            13'h1244: rddata <= 8'h4D;
            13'h1245: rddata <= 8'h20;
            13'h1246: rddata <= 8'hE9;
            13'h1247: rddata <= 8'h29;
            13'h1248: rddata <= 8'h29;
            13'h1249: rddata <= 8'hC1;
            13'h124A: rddata <= 8'h09;
            13'h124B: rddata <= 8'hEB;
            13'h124C: rddata <= 8'h2A;
            13'h124D: rddata <= 8'hD0;
            13'h124E: rddata <= 8'h38;
            13'h124F: rddata <= 8'hC9;
            13'h1250: rddata <= 8'h21;
            13'h1251: rddata <= 8'h57;
            13'h1252: rddata <= 8'h17;
            13'h1253: rddata <= 8'hCD;
            13'h1254: rddata <= 8'h31;
            13'h1255: rddata <= 8'h15;
            13'h1256: rddata <= 8'h18;
            13'h1257: rddata <= 8'h09;
            13'h1258: rddata <= 8'hCD;
            13'h1259: rddata <= 8'h31;
            13'h125A: rddata <= 8'h15;
            13'h125B: rddata <= 8'h21;
            13'h125C: rddata <= 8'hC1;
            13'h125D: rddata <= 8'hD1;
            13'h125E: rddata <= 8'hCD;
            13'h125F: rddata <= 8'h0B;
            13'h1260: rddata <= 8'h15;
            13'h1261: rddata <= 8'h78;
            13'h1262: rddata <= 8'hB7;
            13'h1263: rddata <= 8'hC8;
            13'h1264: rddata <= 8'h3A;
            13'h1265: rddata <= 8'hE7;
            13'h1266: rddata <= 8'h38;
            13'h1267: rddata <= 8'hB7;
            13'h1268: rddata <= 8'hCA;
            13'h1269: rddata <= 8'h23;
            13'h126A: rddata <= 8'h15;
            13'h126B: rddata <= 8'h90;
            13'h126C: rddata <= 8'h30;
            13'h126D: rddata <= 8'h0C;
            13'h126E: rddata <= 8'h2F;
            13'h126F: rddata <= 8'h3C;
            13'h1270: rddata <= 8'hEB;
            13'h1271: rddata <= 8'hCD;
            13'h1272: rddata <= 8'h13;
            13'h1273: rddata <= 8'h15;
            13'h1274: rddata <= 8'hEB;
            13'h1275: rddata <= 8'hCD;
            13'h1276: rddata <= 8'h23;
            13'h1277: rddata <= 8'h15;
            13'h1278: rddata <= 8'hC1;
            13'h1279: rddata <= 8'hD1;
            13'h127A: rddata <= 8'hFE;
            13'h127B: rddata <= 8'h19;
            13'h127C: rddata <= 8'hD0;
            13'h127D: rddata <= 8'hF5;
            13'h127E: rddata <= 8'hCD;
            13'h127F: rddata <= 8'h46;
            13'h1280: rddata <= 8'h15;
            13'h1281: rddata <= 8'h67;
            13'h1282: rddata <= 8'hF1;
            13'h1283: rddata <= 8'hCD;
            13'h1284: rddata <= 8'h30;
            13'h1285: rddata <= 8'h13;
            13'h1286: rddata <= 8'h7C;
            13'h1287: rddata <= 8'hB7;
            13'h1288: rddata <= 8'h21;
            13'h1289: rddata <= 8'hE4;
            13'h128A: rddata <= 8'h38;
            13'h128B: rddata <= 8'hF2;
            13'h128C: rddata <= 8'h9F;
            13'h128D: rddata <= 8'h12;
            13'h128E: rddata <= 8'hCD;
            13'h128F: rddata <= 8'h10;
            13'h1290: rddata <= 8'h13;
            13'h1291: rddata <= 8'h30;
            13'h1292: rddata <= 8'h5E;
            13'h1293: rddata <= 8'h23;
            13'h1294: rddata <= 8'h34;
            13'h1295: rddata <= 8'hCA;
            13'h1296: rddata <= 8'hD3;
            13'h1297: rddata <= 8'h03;
            13'h1298: rddata <= 8'h2E;
            13'h1299: rddata <= 8'h01;
            13'h129A: rddata <= 8'hCD;
            13'h129B: rddata <= 8'h52;
            13'h129C: rddata <= 8'h13;
            13'h129D: rddata <= 8'h18;
            13'h129E: rddata <= 8'h52;
            13'h129F: rddata <= 8'hAF;
            13'h12A0: rddata <= 8'h90;
            13'h12A1: rddata <= 8'h47;
            13'h12A2: rddata <= 8'h7E;
            13'h12A3: rddata <= 8'h9B;
            13'h12A4: rddata <= 8'h5F;
            13'h12A5: rddata <= 8'h23;
            13'h12A6: rddata <= 8'h7E;
            13'h12A7: rddata <= 8'h9A;
            13'h12A8: rddata <= 8'h57;
            13'h12A9: rddata <= 8'h23;
            13'h12AA: rddata <= 8'h7E;
            13'h12AB: rddata <= 8'h99;
            13'h12AC: rddata <= 8'h4F;
            13'h12AD: rddata <= 8'hDC;
            13'h12AE: rddata <= 8'h1C;
            13'h12AF: rddata <= 8'h13;
            13'h12B0: rddata <= 8'h68;
            13'h12B1: rddata <= 8'h63;
            13'h12B2: rddata <= 8'hAF;
            13'h12B3: rddata <= 8'h47;
            13'h12B4: rddata <= 8'h79;
            13'h12B5: rddata <= 8'hB7;
            13'h12B6: rddata <= 8'h20;
            13'h12B7: rddata <= 8'h27;
            13'h12B8: rddata <= 8'h4A;
            13'h12B9: rddata <= 8'h54;
            13'h12BA: rddata <= 8'h65;
            13'h12BB: rddata <= 8'h6F;
            13'h12BC: rddata <= 8'h78;
            13'h12BD: rddata <= 8'hD6;
            13'h12BE: rddata <= 8'h08;
            13'h12BF: rddata <= 8'hFE;
            13'h12C0: rddata <= 8'hE0;
            13'h12C1: rddata <= 8'h20;
            13'h12C2: rddata <= 8'hF0;
            13'h12C3: rddata <= 8'hAF;
            13'h12C4: rddata <= 8'h32;
            13'h12C5: rddata <= 8'hE7;
            13'h12C6: rddata <= 8'h38;
            13'h12C7: rddata <= 8'hC9;
            13'h12C8: rddata <= 8'h7C;
            13'h12C9: rddata <= 8'hB5;
            13'h12CA: rddata <= 8'hB2;
            13'h12CB: rddata <= 8'h20;
            13'h12CC: rddata <= 8'h0A;
            13'h12CD: rddata <= 8'h79;
            13'h12CE: rddata <= 8'h05;
            13'h12CF: rddata <= 8'h17;
            13'h12D0: rddata <= 8'h30;
            13'h12D1: rddata <= 8'hFC;
            13'h12D2: rddata <= 8'h04;
            13'h12D3: rddata <= 8'h1F;
            13'h12D4: rddata <= 8'h4F;
            13'h12D5: rddata <= 8'h18;
            13'h12D6: rddata <= 8'h0B;
            13'h12D7: rddata <= 8'h05;
            13'h12D8: rddata <= 8'h29;
            13'h12D9: rddata <= 8'h7A;
            13'h12DA: rddata <= 8'h17;
            13'h12DB: rddata <= 8'h57;
            13'h12DC: rddata <= 8'h79;
            13'h12DD: rddata <= 8'h8F;
            13'h12DE: rddata <= 8'h4F;
            13'h12DF: rddata <= 8'hF2;
            13'h12E0: rddata <= 8'hC8;
            13'h12E1: rddata <= 8'h12;
            13'h12E2: rddata <= 8'h78;
            13'h12E3: rddata <= 8'h5C;
            13'h12E4: rddata <= 8'h45;
            13'h12E5: rddata <= 8'hB7;
            13'h12E6: rddata <= 8'h28;
            13'h12E7: rddata <= 8'h09;
            13'h12E8: rddata <= 8'h21;
            13'h12E9: rddata <= 8'hE7;
            13'h12EA: rddata <= 8'h38;
            13'h12EB: rddata <= 8'h86;
            13'h12EC: rddata <= 8'h77;
            13'h12ED: rddata <= 8'h30;
            13'h12EE: rddata <= 8'hD4;
            13'h12EF: rddata <= 8'h28;
            13'h12F0: rddata <= 8'hD2;
            13'h12F1: rddata <= 8'h78;
            13'h12F2: rddata <= 8'h21;
            13'h12F3: rddata <= 8'hE7;
            13'h12F4: rddata <= 8'h38;
            13'h12F5: rddata <= 8'hB7;
            13'h12F6: rddata <= 8'hFC;
            13'h12F7: rddata <= 8'h03;
            13'h12F8: rddata <= 8'h13;
            13'h12F9: rddata <= 8'h46;
            13'h12FA: rddata <= 8'h23;
            13'h12FB: rddata <= 8'h7E;
            13'h12FC: rddata <= 8'hE6;
            13'h12FD: rddata <= 8'h80;
            13'h12FE: rddata <= 8'hA9;
            13'h12FF: rddata <= 8'h4F;
            13'h1300: rddata <= 8'hC3;
            13'h1301: rddata <= 8'h23;
            13'h1302: rddata <= 8'h15;
            13'h1303: rddata <= 8'h1C;
            13'h1304: rddata <= 8'hC0;
            13'h1305: rddata <= 8'h14;
            13'h1306: rddata <= 8'hC0;
            13'h1307: rddata <= 8'h0C;
            13'h1308: rddata <= 8'hC0;
            13'h1309: rddata <= 8'h0E;
            13'h130A: rddata <= 8'h80;
            13'h130B: rddata <= 8'h34;
            13'h130C: rddata <= 8'hC0;
            13'h130D: rddata <= 8'hC3;
            13'h130E: rddata <= 8'hD3;
            13'h130F: rddata <= 8'h03;
            13'h1310: rddata <= 8'h7E;
            13'h1311: rddata <= 8'h83;
            13'h1312: rddata <= 8'h5F;
            13'h1313: rddata <= 8'h23;
            13'h1314: rddata <= 8'h7E;
            13'h1315: rddata <= 8'h8A;
            13'h1316: rddata <= 8'h57;
            13'h1317: rddata <= 8'h23;
            13'h1318: rddata <= 8'h7E;
            13'h1319: rddata <= 8'h89;
            13'h131A: rddata <= 8'h4F;
            13'h131B: rddata <= 8'hC9;
            13'h131C: rddata <= 8'h21;
            13'h131D: rddata <= 8'hE8;
            13'h131E: rddata <= 8'h38;
            13'h131F: rddata <= 8'h7E;
            13'h1320: rddata <= 8'h2F;
            13'h1321: rddata <= 8'h77;
            13'h1322: rddata <= 8'hAF;
            13'h1323: rddata <= 8'h6F;
            13'h1324: rddata <= 8'h90;
            13'h1325: rddata <= 8'h47;
            13'h1326: rddata <= 8'h7D;
            13'h1327: rddata <= 8'h9B;
            13'h1328: rddata <= 8'h5F;
            13'h1329: rddata <= 8'h7D;
            13'h132A: rddata <= 8'h9A;
            13'h132B: rddata <= 8'h57;
            13'h132C: rddata <= 8'h7D;
            13'h132D: rddata <= 8'h99;
            13'h132E: rddata <= 8'h4F;
            13'h132F: rddata <= 8'hC9;
            13'h1330: rddata <= 8'h06;
            13'h1331: rddata <= 8'h00;
            13'h1332: rddata <= 8'hD6;
            13'h1333: rddata <= 8'h08;
            13'h1334: rddata <= 8'h38;
            13'h1335: rddata <= 8'h07;
            13'h1336: rddata <= 8'h43;
            13'h1337: rddata <= 8'h5A;
            13'h1338: rddata <= 8'h51;
            13'h1339: rddata <= 8'h0E;
            13'h133A: rddata <= 8'h00;
            13'h133B: rddata <= 8'h18;
            13'h133C: rddata <= 8'hF5;
            13'h133D: rddata <= 8'hC6;
            13'h133E: rddata <= 8'h09;
            13'h133F: rddata <= 8'h6F;
            13'h1340: rddata <= 8'h7A;
            13'h1341: rddata <= 8'hB3;
            13'h1342: rddata <= 8'hB0;
            13'h1343: rddata <= 8'h20;
            13'h1344: rddata <= 8'h09;
            13'h1345: rddata <= 8'h79;
            13'h1346: rddata <= 8'h2D;
            13'h1347: rddata <= 8'hC8;
            13'h1348: rddata <= 8'h1F;
            13'h1349: rddata <= 8'h4F;
            13'h134A: rddata <= 8'h30;
            13'h134B: rddata <= 8'hFA;
            13'h134C: rddata <= 8'h18;
            13'h134D: rddata <= 8'h06;
            13'h134E: rddata <= 8'hAF;
            13'h134F: rddata <= 8'h2D;
            13'h1350: rddata <= 8'hC8;
            13'h1351: rddata <= 8'h79;
            13'h1352: rddata <= 8'h1F;
            13'h1353: rddata <= 8'h4F;
            13'h1354: rddata <= 8'h7A;
            13'h1355: rddata <= 8'h1F;
            13'h1356: rddata <= 8'h57;
            13'h1357: rddata <= 8'h7B;
            13'h1358: rddata <= 8'h1F;
            13'h1359: rddata <= 8'h5F;
            13'h135A: rddata <= 8'h78;
            13'h135B: rddata <= 8'h1F;
            13'h135C: rddata <= 8'h47;
            13'h135D: rddata <= 8'h18;
            13'h135E: rddata <= 8'hEF;
            13'h135F: rddata <= 8'h00;
            13'h1360: rddata <= 8'h00;
            13'h1361: rddata <= 8'h00;
            13'h1362: rddata <= 8'h81;
            13'h1363: rddata <= 8'h04;
            13'h1364: rddata <= 8'h9A;
            13'h1365: rddata <= 8'hF7;
            13'h1366: rddata <= 8'h19;
            13'h1367: rddata <= 8'h83;
            13'h1368: rddata <= 8'h24;
            13'h1369: rddata <= 8'h63;
            13'h136A: rddata <= 8'h43;
            13'h136B: rddata <= 8'h83;
            13'h136C: rddata <= 8'h75;
            13'h136D: rddata <= 8'hCD;
            13'h136E: rddata <= 8'h8D;
            13'h136F: rddata <= 8'h84;
            13'h1370: rddata <= 8'hA9;
            13'h1371: rddata <= 8'h7F;
            13'h1372: rddata <= 8'h83;
            13'h1373: rddata <= 8'h82;
            13'h1374: rddata <= 8'h04;
            13'h1375: rddata <= 8'h00;
            13'h1376: rddata <= 8'h00;
            13'h1377: rddata <= 8'h00;
            13'h1378: rddata <= 8'h81;
            13'h1379: rddata <= 8'hE2;
            13'h137A: rddata <= 8'hB0;
            13'h137B: rddata <= 8'h4D;
            13'h137C: rddata <= 8'h83;
            13'h137D: rddata <= 8'h0A;
            13'h137E: rddata <= 8'h72;
            13'h137F: rddata <= 8'h11;
            13'h1380: rddata <= 8'h83;
            13'h1381: rddata <= 8'hF4;
            13'h1382: rddata <= 8'h04;
            13'h1383: rddata <= 8'h35;
            13'h1384: rddata <= 8'h7F;
            13'h1385: rddata <= 8'hEF;
            13'h1386: rddata <= 8'hB7;
            13'h1387: rddata <= 8'hEA;
            13'h1388: rddata <= 8'h97;
            13'h1389: rddata <= 8'h06;
            13'h138A: rddata <= 8'hCD;
            13'h138B: rddata <= 8'h95;
            13'h138C: rddata <= 8'h13;
            13'h138D: rddata <= 8'h01;
            13'h138E: rddata <= 8'h31;
            13'h138F: rddata <= 8'h80;
            13'h1390: rddata <= 8'h11;
            13'h1391: rddata <= 8'h18;
            13'h1392: rddata <= 8'h72;
            13'h1393: rddata <= 8'h18;
            13'h1394: rddata <= 8'h36;
            13'h1395: rddata <= 8'hCD;
            13'h1396: rddata <= 8'h2E;
            13'h1397: rddata <= 8'h15;
            13'h1398: rddata <= 8'h3E;
            13'h1399: rddata <= 8'h80;
            13'h139A: rddata <= 8'h32;
            13'h139B: rddata <= 8'hE7;
            13'h139C: rddata <= 8'h38;
            13'h139D: rddata <= 8'hA8;
            13'h139E: rddata <= 8'hF5;
            13'h139F: rddata <= 8'hCD;
            13'h13A0: rddata <= 8'h13;
            13'h13A1: rddata <= 8'h15;
            13'h13A2: rddata <= 8'h21;
            13'h13A3: rddata <= 8'h63;
            13'h13A4: rddata <= 8'h13;
            13'h13A5: rddata <= 8'hCD;
            13'h13A6: rddata <= 8'h46;
            13'h13A7: rddata <= 8'h18;
            13'h13A8: rddata <= 8'hC1;
            13'h13A9: rddata <= 8'hE1;
            13'h13AA: rddata <= 8'hCD;
            13'h13AB: rddata <= 8'h13;
            13'h13AC: rddata <= 8'h15;
            13'h13AD: rddata <= 8'hEB;
            13'h13AE: rddata <= 8'hCD;
            13'h13AF: rddata <= 8'h23;
            13'h13B0: rddata <= 8'h15;
            13'h13B1: rddata <= 8'h21;
            13'h13B2: rddata <= 8'h74;
            13'h13B3: rddata <= 8'h13;
            13'h13B4: rddata <= 8'hCD;
            13'h13B5: rddata <= 8'h46;
            13'h13B6: rddata <= 8'h18;
            13'h13B7: rddata <= 8'hC1;
            13'h13B8: rddata <= 8'hD1;
            13'h13B9: rddata <= 8'hCD;
            13'h13BA: rddata <= 8'h2F;
            13'h13BB: rddata <= 8'h14;
            13'h13BC: rddata <= 8'hF1;
            13'h13BD: rddata <= 8'hCD;
            13'h13BE: rddata <= 8'h13;
            13'h13BF: rddata <= 8'h15;
            13'h13C0: rddata <= 8'hCD;
            13'h13C1: rddata <= 8'hF6;
            13'h13C2: rddata <= 8'h14;
            13'h13C3: rddata <= 8'hC1;
            13'h13C4: rddata <= 8'hD1;
            13'h13C5: rddata <= 8'hC3;
            13'h13C6: rddata <= 8'h61;
            13'h13C7: rddata <= 8'h12;
            13'h13C8: rddata <= 8'h21;
            13'h13C9: rddata <= 8'hC1;
            13'h13CA: rddata <= 8'hD1;
            13'h13CB: rddata <= 8'hEF;
            13'h13CC: rddata <= 8'hC8;
            13'h13CD: rddata <= 8'h2E;
            13'h13CE: rddata <= 8'h00;
            13'h13CF: rddata <= 8'hCD;
            13'h13D0: rddata <= 8'hAC;
            13'h13D1: rddata <= 8'h14;
            13'h13D2: rddata <= 8'h79;
            13'h13D3: rddata <= 8'h32;
            13'h13D4: rddata <= 8'hF6;
            13'h13D5: rddata <= 8'h38;
            13'h13D6: rddata <= 8'hEB;
            13'h13D7: rddata <= 8'h22;
            13'h13D8: rddata <= 8'hF7;
            13'h13D9: rddata <= 8'h38;
            13'h13DA: rddata <= 8'h01;
            13'h13DB: rddata <= 8'h00;
            13'h13DC: rddata <= 8'h00;
            13'h13DD: rddata <= 8'h50;
            13'h13DE: rddata <= 8'h58;
            13'h13DF: rddata <= 8'h21;
            13'h13E0: rddata <= 8'hB0;
            13'h13E1: rddata <= 8'h12;
            13'h13E2: rddata <= 8'hE5;
            13'h13E3: rddata <= 8'h21;
            13'h13E4: rddata <= 8'hEB;
            13'h13E5: rddata <= 8'h13;
            13'h13E6: rddata <= 8'hE5;
            13'h13E7: rddata <= 8'hE5;
            13'h13E8: rddata <= 8'h21;
            13'h13E9: rddata <= 8'hE4;
            13'h13EA: rddata <= 8'h38;
            13'h13EB: rddata <= 8'h7E;
            13'h13EC: rddata <= 8'h23;
            13'h13ED: rddata <= 8'hB7;
            13'h13EE: rddata <= 8'h28;
            13'h13EF: rddata <= 8'h2C;
            13'h13F0: rddata <= 8'hE5;
            13'h13F1: rddata <= 8'h2E;
            13'h13F2: rddata <= 8'h08;
            13'h13F3: rddata <= 8'h1F;
            13'h13F4: rddata <= 8'h67;
            13'h13F5: rddata <= 8'h79;
            13'h13F6: rddata <= 8'h30;
            13'h13F7: rddata <= 8'h0B;
            13'h13F8: rddata <= 8'hE5;
            13'h13F9: rddata <= 8'h2A;
            13'h13FA: rddata <= 8'hF7;
            13'h13FB: rddata <= 8'h38;
            13'h13FC: rddata <= 8'h19;
            13'h13FD: rddata <= 8'hEB;
            13'h13FE: rddata <= 8'hE1;
            13'h13FF: rddata <= 8'h3A;
            13'h1400: rddata <= 8'hF6;
            13'h1401: rddata <= 8'h38;
            13'h1402: rddata <= 8'h89;
            13'h1403: rddata <= 8'h1F;
            13'h1404: rddata <= 8'h4F;
            13'h1405: rddata <= 8'h7A;
            13'h1406: rddata <= 8'h1F;
            13'h1407: rddata <= 8'h57;
            13'h1408: rddata <= 8'h7B;
            13'h1409: rddata <= 8'h1F;
            13'h140A: rddata <= 8'h5F;
            13'h140B: rddata <= 8'h78;
            13'h140C: rddata <= 8'h1F;
            13'h140D: rddata <= 8'h47;
            13'h140E: rddata <= 8'hE6;
            13'h140F: rddata <= 8'h10;
            13'h1410: rddata <= 8'h28;
            13'h1411: rddata <= 8'h04;
            13'h1412: rddata <= 8'h78;
            13'h1413: rddata <= 8'hF6;
            13'h1414: rddata <= 8'h20;
            13'h1415: rddata <= 8'h47;
            13'h1416: rddata <= 8'h2D;
            13'h1417: rddata <= 8'h7C;
            13'h1418: rddata <= 8'h20;
            13'h1419: rddata <= 8'hD9;
            13'h141A: rddata <= 8'hE1;
            13'h141B: rddata <= 8'hC9;
            13'h141C: rddata <= 8'h43;
            13'h141D: rddata <= 8'h5A;
            13'h141E: rddata <= 8'h51;
            13'h141F: rddata <= 8'h4F;
            13'h1420: rddata <= 8'hC9;
            13'h1421: rddata <= 8'hCD;
            13'h1422: rddata <= 8'h13;
            13'h1423: rddata <= 8'h15;
            13'h1424: rddata <= 8'h01;
            13'h1425: rddata <= 8'h20;
            13'h1426: rddata <= 8'h84;
            13'h1427: rddata <= 8'h11;
            13'h1428: rddata <= 8'h00;
            13'h1429: rddata <= 8'h00;
            13'h142A: rddata <= 8'hCD;
            13'h142B: rddata <= 8'h23;
            13'h142C: rddata <= 8'h15;
            13'h142D: rddata <= 8'hC1;
            13'h142E: rddata <= 8'hD1;
            13'h142F: rddata <= 8'hEF;
            13'h1430: rddata <= 8'hCA;
            13'h1431: rddata <= 8'hC7;
            13'h1432: rddata <= 8'h03;
            13'h1433: rddata <= 8'h2E;
            13'h1434: rddata <= 8'hFF;
            13'h1435: rddata <= 8'hCD;
            13'h1436: rddata <= 8'hAC;
            13'h1437: rddata <= 8'h14;
            13'h1438: rddata <= 8'h34;
            13'h1439: rddata <= 8'hCA;
            13'h143A: rddata <= 8'hD3;
            13'h143B: rddata <= 8'h03;
            13'h143C: rddata <= 8'h34;
            13'h143D: rddata <= 8'hCA;
            13'h143E: rddata <= 8'hD3;
            13'h143F: rddata <= 8'h03;
            13'h1440: rddata <= 8'h2B;
            13'h1441: rddata <= 8'h7E;
            13'h1442: rddata <= 8'h32;
            13'h1443: rddata <= 8'h19;
            13'h1444: rddata <= 8'h38;
            13'h1445: rddata <= 8'h2B;
            13'h1446: rddata <= 8'h7E;
            13'h1447: rddata <= 8'h32;
            13'h1448: rddata <= 8'h15;
            13'h1449: rddata <= 8'h38;
            13'h144A: rddata <= 8'h2B;
            13'h144B: rddata <= 8'h7E;
            13'h144C: rddata <= 8'h32;
            13'h144D: rddata <= 8'h11;
            13'h144E: rddata <= 8'h38;
            13'h144F: rddata <= 8'h41;
            13'h1450: rddata <= 8'hEB;
            13'h1451: rddata <= 8'hAF;
            13'h1452: rddata <= 8'h4F;
            13'h1453: rddata <= 8'h57;
            13'h1454: rddata <= 8'h5F;
            13'h1455: rddata <= 8'h32;
            13'h1456: rddata <= 8'h1C;
            13'h1457: rddata <= 8'h38;
            13'h1458: rddata <= 8'hE5;
            13'h1459: rddata <= 8'hC5;
            13'h145A: rddata <= 8'h7D;
            13'h145B: rddata <= 8'hCD;
            13'h145C: rddata <= 8'h10;
            13'h145D: rddata <= 8'h38;
            13'h145E: rddata <= 8'hDE;
            13'h145F: rddata <= 8'h00;
            13'h1460: rddata <= 8'h3F;
            13'h1461: rddata <= 8'h30;
            13'h1462: rddata <= 8'h07;
            13'h1463: rddata <= 8'h32;
            13'h1464: rddata <= 8'h1C;
            13'h1465: rddata <= 8'h38;
            13'h1466: rddata <= 8'hF1;
            13'h1467: rddata <= 8'hF1;
            13'h1468: rddata <= 8'h37;
            13'h1469: rddata <= 8'hD2;
            13'h146A: rddata <= 8'hC1;
            13'h146B: rddata <= 8'hE1;
            13'h146C: rddata <= 8'h79;
            13'h146D: rddata <= 8'h3C;
            13'h146E: rddata <= 8'h3D;
            13'h146F: rddata <= 8'h1F;
            13'h1470: rddata <= 8'hF2;
            13'h1471: rddata <= 8'h87;
            13'h1472: rddata <= 8'h14;
            13'h1473: rddata <= 8'h17;
            13'h1474: rddata <= 8'h3A;
            13'h1475: rddata <= 8'h1C;
            13'h1476: rddata <= 8'h38;
            13'h1477: rddata <= 8'h1F;
            13'h1478: rddata <= 8'hE6;
            13'h1479: rddata <= 8'hC0;
            13'h147A: rddata <= 8'hF5;
            13'h147B: rddata <= 8'h78;
            13'h147C: rddata <= 8'hB4;
            13'h147D: rddata <= 8'hB5;
            13'h147E: rddata <= 8'h28;
            13'h147F: rddata <= 8'h02;
            13'h1480: rddata <= 8'h3E;
            13'h1481: rddata <= 8'h20;
            13'h1482: rddata <= 8'hE1;
            13'h1483: rddata <= 8'hB4;
            13'h1484: rddata <= 8'hC3;
            13'h1485: rddata <= 8'hF2;
            13'h1486: rddata <= 8'h12;
            13'h1487: rddata <= 8'h17;
            13'h1488: rddata <= 8'h7B;
            13'h1489: rddata <= 8'h17;
            13'h148A: rddata <= 8'h5F;
            13'h148B: rddata <= 8'h7A;
            13'h148C: rddata <= 8'h17;
            13'h148D: rddata <= 8'h57;
            13'h148E: rddata <= 8'h79;
            13'h148F: rddata <= 8'h17;
            13'h1490: rddata <= 8'h4F;
            13'h1491: rddata <= 8'h29;
            13'h1492: rddata <= 8'h78;
            13'h1493: rddata <= 8'h17;
            13'h1494: rddata <= 8'h47;
            13'h1495: rddata <= 8'h3A;
            13'h1496: rddata <= 8'h1C;
            13'h1497: rddata <= 8'h38;
            13'h1498: rddata <= 8'h17;
            13'h1499: rddata <= 8'h32;
            13'h149A: rddata <= 8'h1C;
            13'h149B: rddata <= 8'h38;
            13'h149C: rddata <= 8'h79;
            13'h149D: rddata <= 8'hB2;
            13'h149E: rddata <= 8'hB3;
            13'h149F: rddata <= 8'h20;
            13'h14A0: rddata <= 8'hB7;
            13'h14A1: rddata <= 8'hE5;
            13'h14A2: rddata <= 8'h21;
            13'h14A3: rddata <= 8'hE7;
            13'h14A4: rddata <= 8'h38;
            13'h14A5: rddata <= 8'h35;
            13'h14A6: rddata <= 8'hE1;
            13'h14A7: rddata <= 8'h20;
            13'h14A8: rddata <= 8'hAF;
            13'h14A9: rddata <= 8'hC3;
            13'h14AA: rddata <= 8'hC3;
            13'h14AB: rddata <= 8'h12;
            13'h14AC: rddata <= 8'h78;
            13'h14AD: rddata <= 8'hB7;
            13'h14AE: rddata <= 8'h28;
            13'h14AF: rddata <= 8'h1D;
            13'h14B0: rddata <= 8'h7D;
            13'h14B1: rddata <= 8'h21;
            13'h14B2: rddata <= 8'hE7;
            13'h14B3: rddata <= 8'h38;
            13'h14B4: rddata <= 8'hAE;
            13'h14B5: rddata <= 8'h80;
            13'h14B6: rddata <= 8'h47;
            13'h14B7: rddata <= 8'h1F;
            13'h14B8: rddata <= 8'hA8;
            13'h14B9: rddata <= 8'h78;
            13'h14BA: rddata <= 8'hF2;
            13'h14BB: rddata <= 8'hCC;
            13'h14BC: rddata <= 8'h14;
            13'h14BD: rddata <= 8'hC6;
            13'h14BE: rddata <= 8'h80;
            13'h14BF: rddata <= 8'h77;
            13'h14C0: rddata <= 8'hCA;
            13'h14C1: rddata <= 8'h1A;
            13'h14C2: rddata <= 8'h14;
            13'h14C3: rddata <= 8'hCD;
            13'h14C4: rddata <= 8'h46;
            13'h14C5: rddata <= 8'h15;
            13'h14C6: rddata <= 8'h77;
            13'h14C7: rddata <= 8'h2B;
            13'h14C8: rddata <= 8'hC9;
            13'h14C9: rddata <= 8'hEF;
            13'h14CA: rddata <= 8'h2F;
            13'h14CB: rddata <= 8'hE1;
            13'h14CC: rddata <= 8'hB7;
            13'h14CD: rddata <= 8'hE1;
            13'h14CE: rddata <= 8'hF2;
            13'h14CF: rddata <= 8'hC3;
            13'h14D0: rddata <= 8'h12;
            13'h14D1: rddata <= 8'hC3;
            13'h14D2: rddata <= 8'hD3;
            13'h14D3: rddata <= 8'h03;
            13'h14D4: rddata <= 8'hCD;
            13'h14D5: rddata <= 8'h2E;
            13'h14D6: rddata <= 8'h15;
            13'h14D7: rddata <= 8'h78;
            13'h14D8: rddata <= 8'hB7;
            13'h14D9: rddata <= 8'hC8;
            13'h14DA: rddata <= 8'hC6;
            13'h14DB: rddata <= 8'h02;
            13'h14DC: rddata <= 8'hDA;
            13'h14DD: rddata <= 8'hD3;
            13'h14DE: rddata <= 8'h03;
            13'h14DF: rddata <= 8'h47;
            13'h14E0: rddata <= 8'hCD;
            13'h14E1: rddata <= 8'h61;
            13'h14E2: rddata <= 8'h12;
            13'h14E3: rddata <= 8'h21;
            13'h14E4: rddata <= 8'hE7;
            13'h14E5: rddata <= 8'h38;
            13'h14E6: rddata <= 8'h34;
            13'h14E7: rddata <= 8'hC0;
            13'h14E8: rddata <= 8'hC3;
            13'h14E9: rddata <= 8'hD3;
            13'h14EA: rddata <= 8'h03;
            13'h14EB: rddata <= 8'h3A;
            13'h14EC: rddata <= 8'hE6;
            13'h14ED: rddata <= 8'h38;
            13'h14EE: rddata <= 8'hFE;
            13'h14EF: rddata <= 8'h2F;
            13'h14F0: rddata <= 8'h17;
            13'h14F1: rddata <= 8'h9F;
            13'h14F2: rddata <= 8'hC0;
            13'h14F3: rddata <= 8'h3C;
            13'h14F4: rddata <= 8'hC9;
            13'h14F5: rddata <= 8'hEF;
            13'h14F6: rddata <= 8'h06;
            13'h14F7: rddata <= 8'h88;
            13'h14F8: rddata <= 8'h11;
            13'h14F9: rddata <= 8'h00;
            13'h14FA: rddata <= 8'h00;
            13'h14FB: rddata <= 8'h21;
            13'h14FC: rddata <= 8'hE7;
            13'h14FD: rddata <= 8'h38;
            13'h14FE: rddata <= 8'h4F;
            13'h14FF: rddata <= 8'h70;
            13'h1500: rddata <= 8'h06;
            13'h1501: rddata <= 8'h00;
            13'h1502: rddata <= 8'h23;
            13'h1503: rddata <= 8'h36;
            13'h1504: rddata <= 8'h80;
            13'h1505: rddata <= 8'h17;
            13'h1506: rddata <= 8'hC3;
            13'h1507: rddata <= 8'hAD;
            13'h1508: rddata <= 8'h12;
            13'h1509: rddata <= 8'hEF;
            13'h150A: rddata <= 8'hF0;
            13'h150B: rddata <= 8'h21;
            13'h150C: rddata <= 8'hE6;
            13'h150D: rddata <= 8'h38;
            13'h150E: rddata <= 8'h7E;
            13'h150F: rddata <= 8'hEE;
            13'h1510: rddata <= 8'h80;
            13'h1511: rddata <= 8'h77;
            13'h1512: rddata <= 8'hC9;
            13'h1513: rddata <= 8'hEB;
            13'h1514: rddata <= 8'h2A;
            13'h1515: rddata <= 8'hE4;
            13'h1516: rddata <= 8'h38;
            13'h1517: rddata <= 8'hE3;
            13'h1518: rddata <= 8'hE5;
            13'h1519: rddata <= 8'h2A;
            13'h151A: rddata <= 8'hE6;
            13'h151B: rddata <= 8'h38;
            13'h151C: rddata <= 8'hE3;
            13'h151D: rddata <= 8'hE5;
            13'h151E: rddata <= 8'hEB;
            13'h151F: rddata <= 8'hC9;
            13'h1520: rddata <= 8'hCD;
            13'h1521: rddata <= 8'h31;
            13'h1522: rddata <= 8'h15;
            13'h1523: rddata <= 8'hEB;
            13'h1524: rddata <= 8'h22;
            13'h1525: rddata <= 8'hE4;
            13'h1526: rddata <= 8'h38;
            13'h1527: rddata <= 8'h60;
            13'h1528: rddata <= 8'h69;
            13'h1529: rddata <= 8'h22;
            13'h152A: rddata <= 8'hE6;
            13'h152B: rddata <= 8'h38;
            13'h152C: rddata <= 8'hEB;
            13'h152D: rddata <= 8'hC9;
            13'h152E: rddata <= 8'h21;
            13'h152F: rddata <= 8'hE4;
            13'h1530: rddata <= 8'h38;
            13'h1531: rddata <= 8'h5E;
            13'h1532: rddata <= 8'h23;
            13'h1533: rddata <= 8'h56;
            13'h1534: rddata <= 8'h23;
            13'h1535: rddata <= 8'h4E;
            13'h1536: rddata <= 8'h23;
            13'h1537: rddata <= 8'h46;
            13'h1538: rddata <= 8'h23;
            13'h1539: rddata <= 8'hC9;
            13'h153A: rddata <= 8'h11;
            13'h153B: rddata <= 8'hE4;
            13'h153C: rddata <= 8'h38;
            13'h153D: rddata <= 8'h06;
            13'h153E: rddata <= 8'h04;
            13'h153F: rddata <= 8'h1A;
            13'h1540: rddata <= 8'h77;
            13'h1541: rddata <= 8'h13;
            13'h1542: rddata <= 8'h23;
            13'h1543: rddata <= 8'h10;
            13'h1544: rddata <= 8'hFA;
            13'h1545: rddata <= 8'hC9;
            13'h1546: rddata <= 8'h21;
            13'h1547: rddata <= 8'hE6;
            13'h1548: rddata <= 8'h38;
            13'h1549: rddata <= 8'h7E;
            13'h154A: rddata <= 8'h07;
            13'h154B: rddata <= 8'h37;
            13'h154C: rddata <= 8'h1F;
            13'h154D: rddata <= 8'h77;
            13'h154E: rddata <= 8'h3F;
            13'h154F: rddata <= 8'h1F;
            13'h1550: rddata <= 8'h23;
            13'h1551: rddata <= 8'h23;
            13'h1552: rddata <= 8'h77;
            13'h1553: rddata <= 8'h79;
            13'h1554: rddata <= 8'h07;
            13'h1555: rddata <= 8'h37;
            13'h1556: rddata <= 8'h1F;
            13'h1557: rddata <= 8'h4F;
            13'h1558: rddata <= 8'h1F;
            13'h1559: rddata <= 8'hAE;
            13'h155A: rddata <= 8'hC9;
            13'h155B: rddata <= 8'h78;
            13'h155C: rddata <= 8'hB7;
            13'h155D: rddata <= 8'hCA;
            13'h155E: rddata <= 8'h28;
            13'h155F: rddata <= 8'h00;
            13'h1560: rddata <= 8'h21;
            13'h1561: rddata <= 8'hEF;
            13'h1562: rddata <= 8'h14;
            13'h1563: rddata <= 8'hE5;
            13'h1564: rddata <= 8'hEF;
            13'h1565: rddata <= 8'h79;
            13'h1566: rddata <= 8'hC8;
            13'h1567: rddata <= 8'h21;
            13'h1568: rddata <= 8'hE6;
            13'h1569: rddata <= 8'h38;
            13'h156A: rddata <= 8'hAE;
            13'h156B: rddata <= 8'h79;
            13'h156C: rddata <= 8'hF8;
            13'h156D: rddata <= 8'hCD;
            13'h156E: rddata <= 8'h73;
            13'h156F: rddata <= 8'h15;
            13'h1570: rddata <= 8'h1F;
            13'h1571: rddata <= 8'hA9;
            13'h1572: rddata <= 8'hC9;
            13'h1573: rddata <= 8'h23;
            13'h1574: rddata <= 8'h78;
            13'h1575: rddata <= 8'hBE;
            13'h1576: rddata <= 8'hC0;
            13'h1577: rddata <= 8'h2B;
            13'h1578: rddata <= 8'h79;
            13'h1579: rddata <= 8'hBE;
            13'h157A: rddata <= 8'hC0;
            13'h157B: rddata <= 8'h2B;
            13'h157C: rddata <= 8'h7A;
            13'h157D: rddata <= 8'hBE;
            13'h157E: rddata <= 8'hC0;
            13'h157F: rddata <= 8'h2B;
            13'h1580: rddata <= 8'h7B;
            13'h1581: rddata <= 8'h96;
            13'h1582: rddata <= 8'hC0;
            13'h1583: rddata <= 8'hE1;
            13'h1584: rddata <= 8'hE1;
            13'h1585: rddata <= 8'hC9;
            13'h1586: rddata <= 8'h47;
            13'h1587: rddata <= 8'h4F;
            13'h1588: rddata <= 8'h57;
            13'h1589: rddata <= 8'h5F;
            13'h158A: rddata <= 8'hB7;
            13'h158B: rddata <= 8'hC8;
            13'h158C: rddata <= 8'hE5;
            13'h158D: rddata <= 8'hCD;
            13'h158E: rddata <= 8'h2E;
            13'h158F: rddata <= 8'h15;
            13'h1590: rddata <= 8'hCD;
            13'h1591: rddata <= 8'h46;
            13'h1592: rddata <= 8'h15;
            13'h1593: rddata <= 8'hAE;
            13'h1594: rddata <= 8'h67;
            13'h1595: rddata <= 8'hFC;
            13'h1596: rddata <= 8'hAA;
            13'h1597: rddata <= 8'h15;
            13'h1598: rddata <= 8'h3E;
            13'h1599: rddata <= 8'h98;
            13'h159A: rddata <= 8'h90;
            13'h159B: rddata <= 8'hCD;
            13'h159C: rddata <= 8'h30;
            13'h159D: rddata <= 8'h13;
            13'h159E: rddata <= 8'h7C;
            13'h159F: rddata <= 8'h17;
            13'h15A0: rddata <= 8'hDC;
            13'h15A1: rddata <= 8'h03;
            13'h15A2: rddata <= 8'h13;
            13'h15A3: rddata <= 8'h06;
            13'h15A4: rddata <= 8'h00;
            13'h15A5: rddata <= 8'hDC;
            13'h15A6: rddata <= 8'h1C;
            13'h15A7: rddata <= 8'h13;
            13'h15A8: rddata <= 8'hE1;
            13'h15A9: rddata <= 8'hC9;
            13'h15AA: rddata <= 8'h1B;
            13'h15AB: rddata <= 8'h7A;
            13'h15AC: rddata <= 8'hA3;
            13'h15AD: rddata <= 8'h3C;
            13'h15AE: rddata <= 8'hC0;
            13'h15AF: rddata <= 8'h0B;
            13'h15B0: rddata <= 8'hC9;
            13'h15B1: rddata <= 8'h21;
            13'h15B2: rddata <= 8'hE7;
            13'h15B3: rddata <= 8'h38;
            13'h15B4: rddata <= 8'h7E;
            13'h15B5: rddata <= 8'hFE;
            13'h15B6: rddata <= 8'h98;
            13'h15B7: rddata <= 8'h3A;
            13'h15B8: rddata <= 8'hE4;
            13'h15B9: rddata <= 8'h38;
            13'h15BA: rddata <= 8'hD0;
            13'h15BB: rddata <= 8'h7E;
            13'h15BC: rddata <= 8'hCD;
            13'h15BD: rddata <= 8'h86;
            13'h15BE: rddata <= 8'h15;
            13'h15BF: rddata <= 8'h36;
            13'h15C0: rddata <= 8'h98;
            13'h15C1: rddata <= 8'h7B;
            13'h15C2: rddata <= 8'hF5;
            13'h15C3: rddata <= 8'h79;
            13'h15C4: rddata <= 8'h17;
            13'h15C5: rddata <= 8'hCD;
            13'h15C6: rddata <= 8'hAD;
            13'h15C7: rddata <= 8'h12;
            13'h15C8: rddata <= 8'hF1;
            13'h15C9: rddata <= 8'hC9;
            13'h15CA: rddata <= 8'h21;
            13'h15CB: rddata <= 8'h00;
            13'h15CC: rddata <= 8'h00;
            13'h15CD: rddata <= 8'h78;
            13'h15CE: rddata <= 8'hB1;
            13'h15CF: rddata <= 8'hC8;
            13'h15D0: rddata <= 8'h3E;
            13'h15D1: rddata <= 8'h10;
            13'h15D2: rddata <= 8'h29;
            13'h15D3: rddata <= 8'hDA;
            13'h15D4: rddata <= 8'hCD;
            13'h15D5: rddata <= 8'h11;
            13'h15D6: rddata <= 8'hEB;
            13'h15D7: rddata <= 8'h29;
            13'h15D8: rddata <= 8'hEB;
            13'h15D9: rddata <= 8'hD2;
            13'h15DA: rddata <= 8'hE0;
            13'h15DB: rddata <= 8'h15;
            13'h15DC: rddata <= 8'h09;
            13'h15DD: rddata <= 8'hDA;
            13'h15DE: rddata <= 8'hCD;
            13'h15DF: rddata <= 8'h11;
            13'h15E0: rddata <= 8'h3D;
            13'h15E1: rddata <= 8'hC2;
            13'h15E2: rddata <= 8'hD2;
            13'h15E3: rddata <= 8'h15;
            13'h15E4: rddata <= 8'hC9;
            13'h15E5: rddata <= 8'hFE;
            13'h15E6: rddata <= 8'h2D;
            13'h15E7: rddata <= 8'hF5;
            13'h15E8: rddata <= 8'h28;
            13'h15E9: rddata <= 8'h05;
            13'h15EA: rddata <= 8'hFE;
            13'h15EB: rddata <= 8'h2B;
            13'h15EC: rddata <= 8'h28;
            13'h15ED: rddata <= 8'h01;
            13'h15EE: rddata <= 8'h2B;
            13'h15EF: rddata <= 8'hCD;
            13'h15F0: rddata <= 8'hC3;
            13'h15F1: rddata <= 8'h12;
            13'h15F2: rddata <= 8'h47;
            13'h15F3: rddata <= 8'h57;
            13'h15F4: rddata <= 8'h5F;
            13'h15F5: rddata <= 8'h2F;
            13'h15F6: rddata <= 8'h4F;
            13'h15F7: rddata <= 8'hD7;
            13'h15F8: rddata <= 8'hDA;
            13'h15F9: rddata <= 8'h3F;
            13'h15FA: rddata <= 8'h16;
            13'h15FB: rddata <= 8'hFE;
            13'h15FC: rddata <= 8'h2E;
            13'h15FD: rddata <= 8'hCA;
            13'h15FE: rddata <= 8'h1A;
            13'h15FF: rddata <= 8'h16;
            13'h1600: rddata <= 8'hFE;
            13'h1601: rddata <= 8'h65;
            13'h1602: rddata <= 8'hCA;
            13'h1603: rddata <= 8'h0A;
            13'h1604: rddata <= 8'h16;
            13'h1605: rddata <= 8'hFE;
            13'h1606: rddata <= 8'h45;
            13'h1607: rddata <= 8'hC2;
            13'h1608: rddata <= 8'h1E;
            13'h1609: rddata <= 8'h16;
            13'h160A: rddata <= 8'hD7;
            13'h160B: rddata <= 8'hCD;
            13'h160C: rddata <= 8'h98;
            13'h160D: rddata <= 8'h0A;
            13'h160E: rddata <= 8'hD7;
            13'h160F: rddata <= 8'hDA;
            13'h1610: rddata <= 8'h61;
            13'h1611: rddata <= 8'h16;
            13'h1612: rddata <= 8'h14;
            13'h1613: rddata <= 8'hC2;
            13'h1614: rddata <= 8'h1E;
            13'h1615: rddata <= 8'h16;
            13'h1616: rddata <= 8'hAF;
            13'h1617: rddata <= 8'h93;
            13'h1618: rddata <= 8'h5F;
            13'h1619: rddata <= 8'h0C;
            13'h161A: rddata <= 8'h0C;
            13'h161B: rddata <= 8'hCA;
            13'h161C: rddata <= 8'hF7;
            13'h161D: rddata <= 8'h15;
            13'h161E: rddata <= 8'hE5;
            13'h161F: rddata <= 8'h7B;
            13'h1620: rddata <= 8'h90;
            13'h1621: rddata <= 8'hF4;
            13'h1622: rddata <= 8'h37;
            13'h1623: rddata <= 8'h16;
            13'h1624: rddata <= 8'hF2;
            13'h1625: rddata <= 8'h2D;
            13'h1626: rddata <= 8'h16;
            13'h1627: rddata <= 8'hF5;
            13'h1628: rddata <= 8'hCD;
            13'h1629: rddata <= 8'h21;
            13'h162A: rddata <= 8'h14;
            13'h162B: rddata <= 8'hF1;
            13'h162C: rddata <= 8'h3C;
            13'h162D: rddata <= 8'hC2;
            13'h162E: rddata <= 8'h21;
            13'h162F: rddata <= 8'h16;
            13'h1630: rddata <= 8'hD1;
            13'h1631: rddata <= 8'hF1;
            13'h1632: rddata <= 8'hCC;
            13'h1633: rddata <= 8'h0B;
            13'h1634: rddata <= 8'h15;
            13'h1635: rddata <= 8'hEB;
            13'h1636: rddata <= 8'hC9;
            13'h1637: rddata <= 8'hC8;
            13'h1638: rddata <= 8'hF5;
            13'h1639: rddata <= 8'hCD;
            13'h163A: rddata <= 8'hD4;
            13'h163B: rddata <= 8'h14;
            13'h163C: rddata <= 8'hF1;
            13'h163D: rddata <= 8'h3D;
            13'h163E: rddata <= 8'hC9;
            13'h163F: rddata <= 8'hD5;
            13'h1640: rddata <= 8'h57;
            13'h1641: rddata <= 8'h78;
            13'h1642: rddata <= 8'h89;
            13'h1643: rddata <= 8'h47;
            13'h1644: rddata <= 8'hC5;
            13'h1645: rddata <= 8'hE5;
            13'h1646: rddata <= 8'hD5;
            13'h1647: rddata <= 8'hCD;
            13'h1648: rddata <= 8'hD4;
            13'h1649: rddata <= 8'h14;
            13'h164A: rddata <= 8'hF1;
            13'h164B: rddata <= 8'hD6;
            13'h164C: rddata <= 8'h30;
            13'h164D: rddata <= 8'hCD;
            13'h164E: rddata <= 8'h56;
            13'h164F: rddata <= 8'h16;
            13'h1650: rddata <= 8'hE1;
            13'h1651: rddata <= 8'hC1;
            13'h1652: rddata <= 8'hD1;
            13'h1653: rddata <= 8'hC3;
            13'h1654: rddata <= 8'hF7;
            13'h1655: rddata <= 8'h15;
            13'h1656: rddata <= 8'hCD;
            13'h1657: rddata <= 8'h13;
            13'h1658: rddata <= 8'h15;
            13'h1659: rddata <= 8'hCD;
            13'h165A: rddata <= 8'hF6;
            13'h165B: rddata <= 8'h14;
            13'h165C: rddata <= 8'hC1;
            13'h165D: rddata <= 8'hD1;
            13'h165E: rddata <= 8'hC3;
            13'h165F: rddata <= 8'h61;
            13'h1660: rddata <= 8'h12;
            13'h1661: rddata <= 8'h7B;
            13'h1662: rddata <= 8'h07;
            13'h1663: rddata <= 8'h07;
            13'h1664: rddata <= 8'h83;
            13'h1665: rddata <= 8'h07;
            13'h1666: rddata <= 8'h86;
            13'h1667: rddata <= 8'hD6;
            13'h1668: rddata <= 8'h30;
            13'h1669: rddata <= 8'h5F;
            13'h166A: rddata <= 8'hC3;
            13'h166B: rddata <= 8'h0E;
            13'h166C: rddata <= 8'h16;
            13'h166D: rddata <= 8'hE5;
            13'h166E: rddata <= 8'h21;
            13'h166F: rddata <= 8'h69;
            13'h1670: rddata <= 8'h03;
            13'h1671: rddata <= 8'hCD;
            13'h1672: rddata <= 8'h9D;
            13'h1673: rddata <= 8'h0E;
            13'h1674: rddata <= 8'hE1;
            13'h1675: rddata <= 8'h11;
            13'h1676: rddata <= 8'h9C;
            13'h1677: rddata <= 8'h0E;
            13'h1678: rddata <= 8'hD5;
            13'h1679: rddata <= 8'hEB;
            13'h167A: rddata <= 8'hAF;
            13'h167B: rddata <= 8'h06;
            13'h167C: rddata <= 8'h98;
            13'h167D: rddata <= 8'hCD;
            13'h167E: rddata <= 8'hFB;
            13'h167F: rddata <= 8'h14;
            13'h1680: rddata <= 8'h21;
            13'h1681: rddata <= 8'hE9;
            13'h1682: rddata <= 8'h38;
            13'h1683: rddata <= 8'hE5;
            13'h1684: rddata <= 8'hEF;
            13'h1685: rddata <= 8'h36;
            13'h1686: rddata <= 8'h20;
            13'h1687: rddata <= 8'hF2;
            13'h1688: rddata <= 8'h8C;
            13'h1689: rddata <= 8'h16;
            13'h168A: rddata <= 8'h36;
            13'h168B: rddata <= 8'h2D;
            13'h168C: rddata <= 8'h23;
            13'h168D: rddata <= 8'h36;
            13'h168E: rddata <= 8'h30;
            13'h168F: rddata <= 8'hCA;
            13'h1690: rddata <= 8'h42;
            13'h1691: rddata <= 8'h17;
            13'h1692: rddata <= 8'hE5;
            13'h1693: rddata <= 8'hFC;
            13'h1694: rddata <= 8'h0B;
            13'h1695: rddata <= 8'h15;
            13'h1696: rddata <= 8'hAF;
            13'h1697: rddata <= 8'hF5;
            13'h1698: rddata <= 8'hCD;
            13'h1699: rddata <= 8'h48;
            13'h169A: rddata <= 8'h17;
            13'h169B: rddata <= 8'h01;
            13'h169C: rddata <= 8'h43;
            13'h169D: rddata <= 8'h91;
            13'h169E: rddata <= 8'h11;
            13'h169F: rddata <= 8'hF8;
            13'h16A0: rddata <= 8'h4F;
            13'h16A1: rddata <= 8'hCD;
            13'h16A2: rddata <= 8'h5B;
            13'h16A3: rddata <= 8'h15;
            13'h16A4: rddata <= 8'hB7;
            13'h16A5: rddata <= 8'hE2;
            13'h16A6: rddata <= 8'hB9;
            13'h16A7: rddata <= 8'h16;
            13'h16A8: rddata <= 8'hF1;
            13'h16A9: rddata <= 8'hCD;
            13'h16AA: rddata <= 8'h38;
            13'h16AB: rddata <= 8'h16;
            13'h16AC: rddata <= 8'hF5;
            13'h16AD: rddata <= 8'hC3;
            13'h16AE: rddata <= 8'h9B;
            13'h16AF: rddata <= 8'h16;
            13'h16B0: rddata <= 8'hCD;
            13'h16B1: rddata <= 8'h21;
            13'h16B2: rddata <= 8'h14;
            13'h16B3: rddata <= 8'hF1;
            13'h16B4: rddata <= 8'h3C;
            13'h16B5: rddata <= 8'hF5;
            13'h16B6: rddata <= 8'hCD;
            13'h16B7: rddata <= 8'h48;
            13'h16B8: rddata <= 8'h17;
            13'h16B9: rddata <= 8'hCD;
            13'h16BA: rddata <= 8'h50;
            13'h16BB: rddata <= 8'h12;
            13'h16BC: rddata <= 8'h3C;
            13'h16BD: rddata <= 8'hCD;
            13'h16BE: rddata <= 8'h86;
            13'h16BF: rddata <= 8'h15;
            13'h16C0: rddata <= 8'hCD;
            13'h16C1: rddata <= 8'h23;
            13'h16C2: rddata <= 8'h15;
            13'h16C3: rddata <= 8'h01;
            13'h16C4: rddata <= 8'h06;
            13'h16C5: rddata <= 8'h03;
            13'h16C6: rddata <= 8'hF1;
            13'h16C7: rddata <= 8'h81;
            13'h16C8: rddata <= 8'h3C;
            13'h16C9: rddata <= 8'hFA;
            13'h16CA: rddata <= 8'hD5;
            13'h16CB: rddata <= 8'h16;
            13'h16CC: rddata <= 8'hFE;
            13'h16CD: rddata <= 8'h08;
            13'h16CE: rddata <= 8'hD2;
            13'h16CF: rddata <= 8'hD5;
            13'h16D0: rddata <= 8'h16;
            13'h16D1: rddata <= 8'h3C;
            13'h16D2: rddata <= 8'h47;
            13'h16D3: rddata <= 8'h3E;
            13'h16D4: rddata <= 8'h02;
            13'h16D5: rddata <= 8'h3D;
            13'h16D6: rddata <= 8'h3D;
            13'h16D7: rddata <= 8'hE1;
            13'h16D8: rddata <= 8'hF5;
            13'h16D9: rddata <= 8'h11;
            13'h16DA: rddata <= 8'h5E;
            13'h16DB: rddata <= 8'h17;
            13'h16DC: rddata <= 8'h05;
            13'h16DD: rddata <= 8'hC2;
            13'h16DE: rddata <= 8'hE6;
            13'h16DF: rddata <= 8'h16;
            13'h16E0: rddata <= 8'h36;
            13'h16E1: rddata <= 8'h2E;
            13'h16E2: rddata <= 8'h23;
            13'h16E3: rddata <= 8'h36;
            13'h16E4: rddata <= 8'h30;
            13'h16E5: rddata <= 8'h23;
            13'h16E6: rddata <= 8'h05;
            13'h16E7: rddata <= 8'h36;
            13'h16E8: rddata <= 8'h2E;
            13'h16E9: rddata <= 8'hCC;
            13'h16EA: rddata <= 8'h38;
            13'h16EB: rddata <= 8'h15;
            13'h16EC: rddata <= 8'hC5;
            13'h16ED: rddata <= 8'hE5;
            13'h16EE: rddata <= 8'hD5;
            13'h16EF: rddata <= 8'hCD;
            13'h16F0: rddata <= 8'h2E;
            13'h16F1: rddata <= 8'h15;
            13'h16F2: rddata <= 8'hE1;
            13'h16F3: rddata <= 8'h06;
            13'h16F4: rddata <= 8'h2F;
            13'h16F5: rddata <= 8'h04;
            13'h16F6: rddata <= 8'h7B;
            13'h16F7: rddata <= 8'h96;
            13'h16F8: rddata <= 8'h5F;
            13'h16F9: rddata <= 8'h23;
            13'h16FA: rddata <= 8'h7A;
            13'h16FB: rddata <= 8'h9E;
            13'h16FC: rddata <= 8'h57;
            13'h16FD: rddata <= 8'h23;
            13'h16FE: rddata <= 8'h79;
            13'h16FF: rddata <= 8'h9E;
            13'h1700: rddata <= 8'h4F;
            13'h1701: rddata <= 8'h2B;
            13'h1702: rddata <= 8'h2B;
            13'h1703: rddata <= 8'hD2;
            13'h1704: rddata <= 8'hF5;
            13'h1705: rddata <= 8'h16;
            13'h1706: rddata <= 8'hCD;
            13'h1707: rddata <= 8'h10;
            13'h1708: rddata <= 8'h13;
            13'h1709: rddata <= 8'h23;
            13'h170A: rddata <= 8'hCD;
            13'h170B: rddata <= 8'h23;
            13'h170C: rddata <= 8'h15;
            13'h170D: rddata <= 8'hEB;
            13'h170E: rddata <= 8'hE1;
            13'h170F: rddata <= 8'h70;
            13'h1710: rddata <= 8'h23;
            13'h1711: rddata <= 8'hC1;
            13'h1712: rddata <= 8'h0D;
            13'h1713: rddata <= 8'hC2;
            13'h1714: rddata <= 8'hE6;
            13'h1715: rddata <= 8'h16;
            13'h1716: rddata <= 8'h05;
            13'h1717: rddata <= 8'hCA;
            13'h1718: rddata <= 8'h26;
            13'h1719: rddata <= 8'h17;
            13'h171A: rddata <= 8'h2B;
            13'h171B: rddata <= 8'h7E;
            13'h171C: rddata <= 8'hFE;
            13'h171D: rddata <= 8'h30;
            13'h171E: rddata <= 8'hCA;
            13'h171F: rddata <= 8'h1A;
            13'h1720: rddata <= 8'h17;
            13'h1721: rddata <= 8'hFE;
            13'h1722: rddata <= 8'h2E;
            13'h1723: rddata <= 8'hC4;
            13'h1724: rddata <= 8'h38;
            13'h1725: rddata <= 8'h15;
            13'h1726: rddata <= 8'hF1;
            13'h1727: rddata <= 8'hCA;
            13'h1728: rddata <= 8'h45;
            13'h1729: rddata <= 8'h17;
            13'h172A: rddata <= 8'h36;
            13'h172B: rddata <= 8'h45;
            13'h172C: rddata <= 8'h23;
            13'h172D: rddata <= 8'h36;
            13'h172E: rddata <= 8'h2B;
            13'h172F: rddata <= 8'hF2;
            13'h1730: rddata <= 8'h36;
            13'h1731: rddata <= 8'h17;
            13'h1732: rddata <= 8'h36;
            13'h1733: rddata <= 8'h2D;
            13'h1734: rddata <= 8'h2F;
            13'h1735: rddata <= 8'h3C;
            13'h1736: rddata <= 8'h06;
            13'h1737: rddata <= 8'h2F;
            13'h1738: rddata <= 8'h04;
            13'h1739: rddata <= 8'hD6;
            13'h173A: rddata <= 8'h0A;
            13'h173B: rddata <= 8'hD2;
            13'h173C: rddata <= 8'h38;
            13'h173D: rddata <= 8'h17;
            13'h173E: rddata <= 8'hC6;
            13'h173F: rddata <= 8'h3A;
            13'h1740: rddata <= 8'h23;
            13'h1741: rddata <= 8'h70;
            13'h1742: rddata <= 8'h23;
            13'h1743: rddata <= 8'h77;
            13'h1744: rddata <= 8'h23;
            13'h1745: rddata <= 8'h71;
            13'h1746: rddata <= 8'hE1;
            13'h1747: rddata <= 8'hC9;
            13'h1748: rddata <= 8'h01;
            13'h1749: rddata <= 8'h74;
            13'h174A: rddata <= 8'h94;
            13'h174B: rddata <= 8'h11;
            13'h174C: rddata <= 8'hF7;
            13'h174D: rddata <= 8'h23;
            13'h174E: rddata <= 8'hCD;
            13'h174F: rddata <= 8'h5B;
            13'h1750: rddata <= 8'h15;
            13'h1751: rddata <= 8'hB7;
            13'h1752: rddata <= 8'hE1;
            13'h1753: rddata <= 8'hE2;
            13'h1754: rddata <= 8'hB0;
            13'h1755: rddata <= 8'h16;
            13'h1756: rddata <= 8'hE9;
            13'h1757: rddata <= 8'h00;
            13'h1758: rddata <= 8'h00;
            13'h1759: rddata <= 8'h00;
            13'h175A: rddata <= 8'h80;
            13'h175B: rddata <= 8'h40;
            13'h175C: rddata <= 8'h42;
            13'h175D: rddata <= 8'h0F;
            13'h175E: rddata <= 8'hA0;
            13'h175F: rddata <= 8'h86;
            13'h1760: rddata <= 8'h01;
            13'h1761: rddata <= 8'h10;
            13'h1762: rddata <= 8'h27;
            13'h1763: rddata <= 8'h00;
            13'h1764: rddata <= 8'hE8;
            13'h1765: rddata <= 8'h03;
            13'h1766: rddata <= 8'h00;
            13'h1767: rddata <= 8'h64;
            13'h1768: rddata <= 8'h00;
            13'h1769: rddata <= 8'h00;
            13'h176A: rddata <= 8'h0A;
            13'h176B: rddata <= 8'h00;
            13'h176C: rddata <= 8'h00;
            13'h176D: rddata <= 8'h01;
            13'h176E: rddata <= 8'h00;
            13'h176F: rddata <= 8'h00;
            13'h1770: rddata <= 8'h21;
            13'h1771: rddata <= 8'h0B;
            13'h1772: rddata <= 8'h15;
            13'h1773: rddata <= 8'hE3;
            13'h1774: rddata <= 8'hE9;
            13'h1775: rddata <= 8'hCD;
            13'h1776: rddata <= 8'h13;
            13'h1777: rddata <= 8'h15;
            13'h1778: rddata <= 8'h21;
            13'h1779: rddata <= 8'h57;
            13'h177A: rddata <= 8'h17;
            13'h177B: rddata <= 8'hCD;
            13'h177C: rddata <= 8'h20;
            13'h177D: rddata <= 8'h15;
            13'h177E: rddata <= 8'hC1;
            13'h177F: rddata <= 8'hD1;
            13'h1780: rddata <= 8'hEF;
            13'h1781: rddata <= 8'h78;
            13'h1782: rddata <= 8'hCA;
            13'h1783: rddata <= 8'hCD;
            13'h1784: rddata <= 8'h17;
            13'h1785: rddata <= 8'hF2;
            13'h1786: rddata <= 8'h8C;
            13'h1787: rddata <= 8'h17;
            13'h1788: rddata <= 8'hB7;
            13'h1789: rddata <= 8'hCA;
            13'h178A: rddata <= 8'hC7;
            13'h178B: rddata <= 8'h03;
            13'h178C: rddata <= 8'hB7;
            13'h178D: rddata <= 8'hCA;
            13'h178E: rddata <= 8'hC4;
            13'h178F: rddata <= 8'h12;
            13'h1790: rddata <= 8'hD5;
            13'h1791: rddata <= 8'hC5;
            13'h1792: rddata <= 8'h79;
            13'h1793: rddata <= 8'hF6;
            13'h1794: rddata <= 8'h7F;
            13'h1795: rddata <= 8'hCD;
            13'h1796: rddata <= 8'h2E;
            13'h1797: rddata <= 8'h15;
            13'h1798: rddata <= 8'hF2;
            13'h1799: rddata <= 8'hB5;
            13'h179A: rddata <= 8'h17;
            13'h179B: rddata <= 8'hF5;
            13'h179C: rddata <= 8'h3A;
            13'h179D: rddata <= 8'hE7;
            13'h179E: rddata <= 8'h38;
            13'h179F: rddata <= 8'hFE;
            13'h17A0: rddata <= 8'h99;
            13'h17A1: rddata <= 8'h38;
            13'h17A2: rddata <= 8'h03;
            13'h17A3: rddata <= 8'hF1;
            13'h17A4: rddata <= 8'h18;
            13'h17A5: rddata <= 8'h0F;
            13'h17A6: rddata <= 8'hF1;
            13'h17A7: rddata <= 8'hD5;
            13'h17A8: rddata <= 8'hC5;
            13'h17A9: rddata <= 8'hCD;
            13'h17AA: rddata <= 8'hB1;
            13'h17AB: rddata <= 8'h15;
            13'h17AC: rddata <= 8'hC1;
            13'h17AD: rddata <= 8'hD1;
            13'h17AE: rddata <= 8'hF5;
            13'h17AF: rddata <= 8'hCD;
            13'h17B0: rddata <= 8'h5B;
            13'h17B1: rddata <= 8'h15;
            13'h17B2: rddata <= 8'hE1;
            13'h17B3: rddata <= 8'h7C;
            13'h17B4: rddata <= 8'h1F;
            13'h17B5: rddata <= 8'hE1;
            13'h17B6: rddata <= 8'h22;
            13'h17B7: rddata <= 8'hE6;
            13'h17B8: rddata <= 8'h38;
            13'h17B9: rddata <= 8'hE1;
            13'h17BA: rddata <= 8'h22;
            13'h17BB: rddata <= 8'hE4;
            13'h17BC: rddata <= 8'h38;
            13'h17BD: rddata <= 8'hDC;
            13'h17BE: rddata <= 8'h70;
            13'h17BF: rddata <= 8'h17;
            13'h17C0: rddata <= 8'hCC;
            13'h17C1: rddata <= 8'h0B;
            13'h17C2: rddata <= 8'h15;
            13'h17C3: rddata <= 8'hD5;
            13'h17C4: rddata <= 8'hC5;
            13'h17C5: rddata <= 8'hCD;
            13'h17C6: rddata <= 8'h85;
            13'h17C7: rddata <= 8'h13;
            13'h17C8: rddata <= 8'hC1;
            13'h17C9: rddata <= 8'hD1;
            13'h17CA: rddata <= 8'hCD;
            13'h17CB: rddata <= 8'hCB;
            13'h17CC: rddata <= 8'h13;
            13'h17CD: rddata <= 8'h01;
            13'h17CE: rddata <= 8'h38;
            13'h17CF: rddata <= 8'h81;
            13'h17D0: rddata <= 8'h11;
            13'h17D1: rddata <= 8'h3B;
            13'h17D2: rddata <= 8'hAA;
            13'h17D3: rddata <= 8'hCD;
            13'h17D4: rddata <= 8'hCB;
            13'h17D5: rddata <= 8'h13;
            13'h17D6: rddata <= 8'h3A;
            13'h17D7: rddata <= 8'hE7;
            13'h17D8: rddata <= 8'h38;
            13'h17D9: rddata <= 8'hFE;
            13'h17DA: rddata <= 8'h88;
            13'h17DB: rddata <= 8'h30;
            13'h17DC: rddata <= 8'h22;
            13'h17DD: rddata <= 8'hFE;
            13'h17DE: rddata <= 8'h68;
            13'h17DF: rddata <= 8'h38;
            13'h17E0: rddata <= 8'h30;
            13'h17E1: rddata <= 8'hCD;
            13'h17E2: rddata <= 8'h13;
            13'h17E3: rddata <= 8'h15;
            13'h17E4: rddata <= 8'hCD;
            13'h17E5: rddata <= 8'hB1;
            13'h17E6: rddata <= 8'h15;
            13'h17E7: rddata <= 8'hC6;
            13'h17E8: rddata <= 8'h81;
            13'h17E9: rddata <= 8'hC1;
            13'h17EA: rddata <= 8'hD1;
            13'h17EB: rddata <= 8'h28;
            13'h17EC: rddata <= 8'h15;
            13'h17ED: rddata <= 8'hF5;
            13'h17EE: rddata <= 8'hCD;
            13'h17EF: rddata <= 8'h5E;
            13'h17F0: rddata <= 8'h12;
            13'h17F1: rddata <= 8'h21;
            13'h17F2: rddata <= 8'h1A;
            13'h17F3: rddata <= 8'h18;
            13'h17F4: rddata <= 8'hCD;
            13'h17F5: rddata <= 8'h46;
            13'h17F6: rddata <= 8'h18;
            13'h17F7: rddata <= 8'hC1;
            13'h17F8: rddata <= 8'h11;
            13'h17F9: rddata <= 8'h00;
            13'h17FA: rddata <= 8'h00;
            13'h17FB: rddata <= 8'h4A;
            13'h17FC: rddata <= 8'hC3;
            13'h17FD: rddata <= 8'hCB;
            13'h17FE: rddata <= 8'h13;
            13'h17FF: rddata <= 8'hCD;
            13'h1800: rddata <= 8'h13;
            13'h1801: rddata <= 8'h15;
            13'h1802: rddata <= 8'h3A;
            13'h1803: rddata <= 8'hE6;
            13'h1804: rddata <= 8'h38;
            13'h1805: rddata <= 8'hB7;
            13'h1806: rddata <= 8'hF2;
            13'h1807: rddata <= 8'h0E;
            13'h1808: rddata <= 8'h18;
            13'h1809: rddata <= 8'hF1;
            13'h180A: rddata <= 8'hF1;
            13'h180B: rddata <= 8'hC3;
            13'h180C: rddata <= 8'hC3;
            13'h180D: rddata <= 8'h12;
            13'h180E: rddata <= 8'hC3;
            13'h180F: rddata <= 8'hD3;
            13'h1810: rddata <= 8'h03;
            13'h1811: rddata <= 8'h01;
            13'h1812: rddata <= 8'h00;
            13'h1813: rddata <= 8'h81;
            13'h1814: rddata <= 8'h11;
            13'h1815: rddata <= 8'h00;
            13'h1816: rddata <= 8'h00;
            13'h1817: rddata <= 8'hC3;
            13'h1818: rddata <= 8'h23;
            13'h1819: rddata <= 8'h15;
            13'h181A: rddata <= 8'h07;
            13'h181B: rddata <= 8'h7C;
            13'h181C: rddata <= 8'h88;
            13'h181D: rddata <= 8'h59;
            13'h181E: rddata <= 8'h74;
            13'h181F: rddata <= 8'hE0;
            13'h1820: rddata <= 8'h97;
            13'h1821: rddata <= 8'h26;
            13'h1822: rddata <= 8'h77;
            13'h1823: rddata <= 8'hC4;
            13'h1824: rddata <= 8'h1D;
            13'h1825: rddata <= 8'h1E;
            13'h1826: rddata <= 8'h7A;
            13'h1827: rddata <= 8'h5E;
            13'h1828: rddata <= 8'h50;
            13'h1829: rddata <= 8'h63;
            13'h182A: rddata <= 8'h7C;
            13'h182B: rddata <= 8'h1A;
            13'h182C: rddata <= 8'hFE;
            13'h182D: rddata <= 8'h75;
            13'h182E: rddata <= 8'h7E;
            13'h182F: rddata <= 8'h18;
            13'h1830: rddata <= 8'h72;
            13'h1831: rddata <= 8'h31;
            13'h1832: rddata <= 8'h80;
            13'h1833: rddata <= 8'h00;
            13'h1834: rddata <= 8'h00;
            13'h1835: rddata <= 8'h00;
            13'h1836: rddata <= 8'h81;
            13'h1837: rddata <= 8'hCD;
            13'h1838: rddata <= 8'h13;
            13'h1839: rddata <= 8'h15;
            13'h183A: rddata <= 8'h11;
            13'h183B: rddata <= 8'hC9;
            13'h183C: rddata <= 8'h13;
            13'h183D: rddata <= 8'hD5;
            13'h183E: rddata <= 8'hE5;
            13'h183F: rddata <= 8'hCD;
            13'h1840: rddata <= 8'h2E;
            13'h1841: rddata <= 8'h15;
            13'h1842: rddata <= 8'hCD;
            13'h1843: rddata <= 8'hCB;
            13'h1844: rddata <= 8'h13;
            13'h1845: rddata <= 8'hE1;
            13'h1846: rddata <= 8'hCD;
            13'h1847: rddata <= 8'h13;
            13'h1848: rddata <= 8'h15;
            13'h1849: rddata <= 8'h7E;
            13'h184A: rddata <= 8'h23;
            13'h184B: rddata <= 8'hCD;
            13'h184C: rddata <= 8'h20;
            13'h184D: rddata <= 8'h15;
            13'h184E: rddata <= 8'h06;
            13'h184F: rddata <= 8'hF1;
            13'h1850: rddata <= 8'hC1;
            13'h1851: rddata <= 8'hD1;
            13'h1852: rddata <= 8'h3D;
            13'h1853: rddata <= 8'hC8;
            13'h1854: rddata <= 8'hD5;
            13'h1855: rddata <= 8'hC5;
            13'h1856: rddata <= 8'hF5;
            13'h1857: rddata <= 8'hE5;
            13'h1858: rddata <= 8'hCD;
            13'h1859: rddata <= 8'hCB;
            13'h185A: rddata <= 8'h13;
            13'h185B: rddata <= 8'hE1;
            13'h185C: rddata <= 8'hCD;
            13'h185D: rddata <= 8'h31;
            13'h185E: rddata <= 8'h15;
            13'h185F: rddata <= 8'hE5;
            13'h1860: rddata <= 8'hCD;
            13'h1861: rddata <= 8'h61;
            13'h1862: rddata <= 8'h12;
            13'h1863: rddata <= 8'hE1;
            13'h1864: rddata <= 8'h18;
            13'h1865: rddata <= 8'hE9;
            13'h1866: rddata <= 8'hEF;
            13'h1867: rddata <= 8'h21;
            13'h1868: rddata <= 8'h20;
            13'h1869: rddata <= 8'h38;
            13'h186A: rddata <= 8'hFA;
            13'h186B: rddata <= 8'hC4;
            13'h186C: rddata <= 8'h18;
            13'h186D: rddata <= 8'h21;
            13'h186E: rddata <= 8'h41;
            13'h186F: rddata <= 8'h38;
            13'h1870: rddata <= 8'hCD;
            13'h1871: rddata <= 8'h20;
            13'h1872: rddata <= 8'h15;
            13'h1873: rddata <= 8'h21;
            13'h1874: rddata <= 8'h20;
            13'h1875: rddata <= 8'h38;
            13'h1876: rddata <= 8'hC8;
            13'h1877: rddata <= 8'h86;
            13'h1878: rddata <= 8'hE6;
            13'h1879: rddata <= 8'h07;
            13'h187A: rddata <= 8'h06;
            13'h187B: rddata <= 8'h00;
            13'h187C: rddata <= 8'h77;
            13'h187D: rddata <= 8'h23;
            13'h187E: rddata <= 8'h87;
            13'h187F: rddata <= 8'h87;
            13'h1880: rddata <= 8'h4F;
            13'h1881: rddata <= 8'h09;
            13'h1882: rddata <= 8'hCD;
            13'h1883: rddata <= 8'h31;
            13'h1884: rddata <= 8'h15;
            13'h1885: rddata <= 8'hCD;
            13'h1886: rddata <= 8'hCB;
            13'h1887: rddata <= 8'h13;
            13'h1888: rddata <= 8'h3A;
            13'h1889: rddata <= 8'h1F;
            13'h188A: rddata <= 8'h38;
            13'h188B: rddata <= 8'h3C;
            13'h188C: rddata <= 8'hE6;
            13'h188D: rddata <= 8'h03;
            13'h188E: rddata <= 8'h06;
            13'h188F: rddata <= 8'h00;
            13'h1890: rddata <= 8'hFE;
            13'h1891: rddata <= 8'h01;
            13'h1892: rddata <= 8'h88;
            13'h1893: rddata <= 8'h32;
            13'h1894: rddata <= 8'h1F;
            13'h1895: rddata <= 8'h38;
            13'h1896: rddata <= 8'h21;
            13'h1897: rddata <= 8'hC7;
            13'h1898: rddata <= 8'h18;
            13'h1899: rddata <= 8'h87;
            13'h189A: rddata <= 8'h87;
            13'h189B: rddata <= 8'h4F;
            13'h189C: rddata <= 8'h09;
            13'h189D: rddata <= 8'hCD;
            13'h189E: rddata <= 8'h53;
            13'h189F: rddata <= 8'h12;
            13'h18A0: rddata <= 8'hCD;
            13'h18A1: rddata <= 8'h2E;
            13'h18A2: rddata <= 8'h15;
            13'h18A3: rddata <= 8'h7B;
            13'h18A4: rddata <= 8'h59;
            13'h18A5: rddata <= 8'hEE;
            13'h18A6: rddata <= 8'h4F;
            13'h18A7: rddata <= 8'h4F;
            13'h18A8: rddata <= 8'h36;
            13'h18A9: rddata <= 8'h80;
            13'h18AA: rddata <= 8'h2B;
            13'h18AB: rddata <= 8'h46;
            13'h18AC: rddata <= 8'h36;
            13'h18AD: rddata <= 8'h80;
            13'h18AE: rddata <= 8'h21;
            13'h18AF: rddata <= 8'h1E;
            13'h18B0: rddata <= 8'h38;
            13'h18B1: rddata <= 8'h34;
            13'h18B2: rddata <= 8'h7E;
            13'h18B3: rddata <= 8'hD6;
            13'h18B4: rddata <= 8'hAB;
            13'h18B5: rddata <= 8'h20;
            13'h18B6: rddata <= 8'h04;
            13'h18B7: rddata <= 8'h77;
            13'h18B8: rddata <= 8'h0C;
            13'h18B9: rddata <= 8'h15;
            13'h18BA: rddata <= 8'h1C;
            13'h18BB: rddata <= 8'hCD;
            13'h18BC: rddata <= 8'hB0;
            13'h18BD: rddata <= 8'h12;
            13'h18BE: rddata <= 8'h21;
            13'h18BF: rddata <= 8'h41;
            13'h18C0: rddata <= 8'h38;
            13'h18C1: rddata <= 8'hC3;
            13'h18C2: rddata <= 8'h3A;
            13'h18C3: rddata <= 8'h15;
            13'h18C4: rddata <= 8'h77;
            13'h18C5: rddata <= 8'h2B;
            13'h18C6: rddata <= 8'h77;
            13'h18C7: rddata <= 8'h2B;
            13'h18C8: rddata <= 8'h77;
            13'h18C9: rddata <= 8'h18;
            13'h18CA: rddata <= 8'hD5;
            13'h18CB: rddata <= 8'h68;
            13'h18CC: rddata <= 8'hB1;
            13'h18CD: rddata <= 8'h46;
            13'h18CE: rddata <= 8'h68;
            13'h18CF: rddata <= 8'h99;
            13'h18D0: rddata <= 8'hE9;
            13'h18D1: rddata <= 8'h92;
            13'h18D2: rddata <= 8'h69;
            13'h18D3: rddata <= 8'h10;
            13'h18D4: rddata <= 8'hD1;
            13'h18D5: rddata <= 8'h75;
            13'h18D6: rddata <= 8'h68;
            13'h18D7: rddata <= 8'h21;
            13'h18D8: rddata <= 8'h53;
            13'h18D9: rddata <= 8'h19;
            13'h18DA: rddata <= 8'hCD;
            13'h18DB: rddata <= 8'h53;
            13'h18DC: rddata <= 8'h12;
            13'h18DD: rddata <= 8'h3A;
            13'h18DE: rddata <= 8'hE7;
            13'h18DF: rddata <= 8'h38;
            13'h18E0: rddata <= 8'hFE;
            13'h18E1: rddata <= 8'h77;
            13'h18E2: rddata <= 8'hD8;
            13'h18E3: rddata <= 8'h3A;
            13'h18E4: rddata <= 8'hE6;
            13'h18E5: rddata <= 8'h38;
            13'h18E6: rddata <= 8'hB7;
            13'h18E7: rddata <= 8'hF2;
            13'h18E8: rddata <= 8'hF3;
            13'h18E9: rddata <= 8'h18;
            13'h18EA: rddata <= 8'hE6;
            13'h18EB: rddata <= 8'h7F;
            13'h18EC: rddata <= 8'h32;
            13'h18ED: rddata <= 8'hE6;
            13'h18EE: rddata <= 8'h38;
            13'h18EF: rddata <= 8'h11;
            13'h18F0: rddata <= 8'h0B;
            13'h18F1: rddata <= 8'h15;
            13'h18F2: rddata <= 8'hD5;
            13'h18F3: rddata <= 8'h01;
            13'h18F4: rddata <= 8'h22;
            13'h18F5: rddata <= 8'h7E;
            13'h18F6: rddata <= 8'h11;
            13'h18F7: rddata <= 8'h83;
            13'h18F8: rddata <= 8'hF9;
            13'h18F9: rddata <= 8'hCD;
            13'h18FA: rddata <= 8'hCB;
            13'h18FB: rddata <= 8'h13;
            13'h18FC: rddata <= 8'hCD;
            13'h18FD: rddata <= 8'h13;
            13'h18FE: rddata <= 8'h15;
            13'h18FF: rddata <= 8'hCD;
            13'h1900: rddata <= 8'hB1;
            13'h1901: rddata <= 8'h15;
            13'h1902: rddata <= 8'hC1;
            13'h1903: rddata <= 8'hD1;
            13'h1904: rddata <= 8'hCD;
            13'h1905: rddata <= 8'h5E;
            13'h1906: rddata <= 8'h12;
            13'h1907: rddata <= 8'h01;
            13'h1908: rddata <= 8'h00;
            13'h1909: rddata <= 8'h7F;
            13'h190A: rddata <= 8'h11;
            13'h190B: rddata <= 8'h00;
            13'h190C: rddata <= 8'h00;
            13'h190D: rddata <= 8'hCD;
            13'h190E: rddata <= 8'h5B;
            13'h190F: rddata <= 8'h15;
            13'h1910: rddata <= 8'hFA;
            13'h1911: rddata <= 8'h35;
            13'h1912: rddata <= 8'h19;
            13'h1913: rddata <= 8'h01;
            13'h1914: rddata <= 8'h80;
            13'h1915: rddata <= 8'h7F;
            13'h1916: rddata <= 8'h11;
            13'h1917: rddata <= 8'h00;
            13'h1918: rddata <= 8'h00;
            13'h1919: rddata <= 8'hCD;
            13'h191A: rddata <= 8'h61;
            13'h191B: rddata <= 8'h12;
            13'h191C: rddata <= 8'h01;
            13'h191D: rddata <= 8'h80;
            13'h191E: rddata <= 8'h80;
            13'h191F: rddata <= 8'h11;
            13'h1920: rddata <= 8'h00;
            13'h1921: rddata <= 8'h00;
            13'h1922: rddata <= 8'hCD;
            13'h1923: rddata <= 8'h61;
            13'h1924: rddata <= 8'h12;
            13'h1925: rddata <= 8'hEF;
            13'h1926: rddata <= 8'hF4;
            13'h1927: rddata <= 8'h0B;
            13'h1928: rddata <= 8'h15;
            13'h1929: rddata <= 8'h01;
            13'h192A: rddata <= 8'h00;
            13'h192B: rddata <= 8'h7F;
            13'h192C: rddata <= 8'h11;
            13'h192D: rddata <= 8'h00;
            13'h192E: rddata <= 8'h00;
            13'h192F: rddata <= 8'hCD;
            13'h1930: rddata <= 8'h61;
            13'h1931: rddata <= 8'h12;
            13'h1932: rddata <= 8'hCD;
            13'h1933: rddata <= 8'h0B;
            13'h1934: rddata <= 8'h15;
            13'h1935: rddata <= 8'h3A;
            13'h1936: rddata <= 8'hE6;
            13'h1937: rddata <= 8'h38;
            13'h1938: rddata <= 8'hB7;
            13'h1939: rddata <= 8'hF5;
            13'h193A: rddata <= 8'hF2;
            13'h193B: rddata <= 8'h42;
            13'h193C: rddata <= 8'h19;
            13'h193D: rddata <= 8'hEE;
            13'h193E: rddata <= 8'h80;
            13'h193F: rddata <= 8'h32;
            13'h1940: rddata <= 8'hE6;
            13'h1941: rddata <= 8'h38;
            13'h1942: rddata <= 8'h21;
            13'h1943: rddata <= 8'h5B;
            13'h1944: rddata <= 8'h19;
            13'h1945: rddata <= 8'hCD;
            13'h1946: rddata <= 8'h37;
            13'h1947: rddata <= 8'h18;
            13'h1948: rddata <= 8'hF1;
            13'h1949: rddata <= 8'hF0;
            13'h194A: rddata <= 8'h3A;
            13'h194B: rddata <= 8'hE6;
            13'h194C: rddata <= 8'h38;
            13'h194D: rddata <= 8'hEE;
            13'h194E: rddata <= 8'h80;
            13'h194F: rddata <= 8'h32;
            13'h1950: rddata <= 8'hE6;
            13'h1951: rddata <= 8'h38;
            13'h1952: rddata <= 8'hC9;
            13'h1953: rddata <= 8'hDB;
            13'h1954: rddata <= 8'h0F;
            13'h1955: rddata <= 8'h49;
            13'h1956: rddata <= 8'h81;
            13'h1957: rddata <= 8'h00;
            13'h1958: rddata <= 8'h00;
            13'h1959: rddata <= 8'h00;
            13'h195A: rddata <= 8'h7F;
            13'h195B: rddata <= 8'h05;
            13'h195C: rddata <= 8'hFB;
            13'h195D: rddata <= 8'hD7;
            13'h195E: rddata <= 8'h1E;
            13'h195F: rddata <= 8'h86;
            13'h1960: rddata <= 8'h65;
            13'h1961: rddata <= 8'h26;
            13'h1962: rddata <= 8'h99;
            13'h1963: rddata <= 8'h87;
            13'h1964: rddata <= 8'h58;
            13'h1965: rddata <= 8'h34;
            13'h1966: rddata <= 8'h23;
            13'h1967: rddata <= 8'h87;
            13'h1968: rddata <= 8'hE1;
            13'h1969: rddata <= 8'h5D;
            13'h196A: rddata <= 8'hA5;
            13'h196B: rddata <= 8'h86;
            13'h196C: rddata <= 8'hDB;
            13'h196D: rddata <= 8'h0F;
            13'h196E: rddata <= 8'h49;
            13'h196F: rddata <= 8'h83;
            13'h1970: rddata <= 8'hCD;
            13'h1971: rddata <= 8'h13;
            13'h1972: rddata <= 8'h15;
            13'h1973: rddata <= 8'hCD;
            13'h1974: rddata <= 8'hDD;
            13'h1975: rddata <= 8'h18;
            13'h1976: rddata <= 8'hC1;
            13'h1977: rddata <= 8'hE1;
            13'h1978: rddata <= 8'hCD;
            13'h1979: rddata <= 8'h13;
            13'h197A: rddata <= 8'h15;
            13'h197B: rddata <= 8'hEB;
            13'h197C: rddata <= 8'hCD;
            13'h197D: rddata <= 8'h23;
            13'h197E: rddata <= 8'h15;
            13'h197F: rddata <= 8'hCD;
            13'h1980: rddata <= 8'hD7;
            13'h1981: rddata <= 8'h18;
            13'h1982: rddata <= 8'hC3;
            13'h1983: rddata <= 8'h2D;
            13'h1984: rddata <= 8'h14;
            13'h1985: rddata <= 8'hF7;
            13'h1986: rddata <= 8'h0E;
            13'h1987: rddata <= 8'hC3;
            13'h1988: rddata <= 8'hC4;
            13'h1989: rddata <= 8'h03;
            13'h198A: rddata <= 8'hF7;
            13'h198B: rddata <= 8'h0D;
            13'h198C: rddata <= 8'hF5;
            13'h198D: rddata <= 8'h3A;
            13'h198E: rddata <= 8'h47;
            13'h198F: rddata <= 8'h38;
            13'h1990: rddata <= 8'hB7;
            13'h1991: rddata <= 8'hCA;
            13'h1992: rddata <= 8'hD6;
            13'h1993: rddata <= 8'h19;
            13'h1994: rddata <= 8'hF1;
            13'h1995: rddata <= 8'hF5;
            13'h1996: rddata <= 8'hFE;
            13'h1997: rddata <= 8'h09;
            13'h1998: rddata <= 8'h20;
            13'h1999: rddata <= 8'h0C;
            13'h199A: rddata <= 8'h3E;
            13'h199B: rddata <= 8'h20;
            13'h199C: rddata <= 8'hDF;
            13'h199D: rddata <= 8'h3A;
            13'h199E: rddata <= 8'h46;
            13'h199F: rddata <= 8'h38;
            13'h19A0: rddata <= 8'hE6;
            13'h19A1: rddata <= 8'h07;
            13'h19A2: rddata <= 8'h20;
            13'h19A3: rddata <= 8'hF6;
            13'h19A4: rddata <= 8'hF1;
            13'h19A5: rddata <= 8'hC9;
            13'h19A6: rddata <= 8'hF1;
            13'h19A7: rddata <= 8'hF5;
            13'h19A8: rddata <= 8'hD6;
            13'h19A9: rddata <= 8'h0D;
            13'h19AA: rddata <= 8'h28;
            13'h19AB: rddata <= 8'h0B;
            13'h19AC: rddata <= 8'h38;
            13'h19AD: rddata <= 8'h0C;
            13'h19AE: rddata <= 8'h3A;
            13'h19AF: rddata <= 8'h46;
            13'h19B0: rddata <= 8'h38;
            13'h19B1: rddata <= 8'h3C;
            13'h19B2: rddata <= 8'hFE;
            13'h19B3: rddata <= 8'h84;
            13'h19B4: rddata <= 8'hCC;
            13'h19B5: rddata <= 8'hC7;
            13'h19B6: rddata <= 8'h19;
            13'h19B7: rddata <= 8'h32;
            13'h19B8: rddata <= 8'h46;
            13'h19B9: rddata <= 8'h38;
            13'h19BA: rddata <= 8'hF1;
            13'h19BB: rddata <= 8'hC3;
            13'h19BC: rddata <= 8'hE8;
            13'h19BD: rddata <= 8'h1A;
            13'h19BE: rddata <= 8'hAF;
            13'h19BF: rddata <= 8'h32;
            13'h19C0: rddata <= 8'h47;
            13'h19C1: rddata <= 8'h38;
            13'h19C2: rddata <= 8'h3A;
            13'h19C3: rddata <= 8'h46;
            13'h19C4: rddata <= 8'h38;
            13'h19C5: rddata <= 8'hB7;
            13'h19C6: rddata <= 8'hC8;
            13'h19C7: rddata <= 8'h3E;
            13'h19C8: rddata <= 8'h0D;
            13'h19C9: rddata <= 8'hCD;
            13'h19CA: rddata <= 8'hBB;
            13'h19CB: rddata <= 8'h19;
            13'h19CC: rddata <= 8'h3E;
            13'h19CD: rddata <= 8'h0A;
            13'h19CE: rddata <= 8'hCD;
            13'h19CF: rddata <= 8'hBB;
            13'h19D0: rddata <= 8'h19;
            13'h19D1: rddata <= 8'hAF;
            13'h19D2: rddata <= 8'h32;
            13'h19D3: rddata <= 8'h46;
            13'h19D4: rddata <= 8'h38;
            13'h19D5: rddata <= 8'hC9;
            13'h19D6: rddata <= 8'hF1;
            13'h19D7: rddata <= 8'hC3;
            13'h19D8: rddata <= 8'h72;
            13'h19D9: rddata <= 8'h1D;
            13'h19DA: rddata <= 8'hCD;
            13'h19DB: rddata <= 8'h2F;
            13'h19DC: rddata <= 8'h1A;
            13'h19DD: rddata <= 8'hC9;
            13'h19DE: rddata <= 8'h3A;
            13'h19DF: rddata <= 8'h00;
            13'h19E0: rddata <= 8'h38;
            13'h19E1: rddata <= 8'hB7;
            13'h19E2: rddata <= 8'hC8;
            13'h19E3: rddata <= 8'h18;
            13'h19E4: rddata <= 8'h05;
            13'h19E5: rddata <= 8'h36;
            13'h19E6: rddata <= 8'h00;
            13'h19E7: rddata <= 8'h21;
            13'h19E8: rddata <= 8'h5F;
            13'h19E9: rddata <= 8'h38;
            13'h19EA: rddata <= 8'h3E;
            13'h19EB: rddata <= 8'h0D;
            13'h19EC: rddata <= 8'hDF;
            13'h19ED: rddata <= 8'h3E;
            13'h19EE: rddata <= 8'h0A;
            13'h19EF: rddata <= 8'hDF;
            13'h19F0: rddata <= 8'h3A;
            13'h19F1: rddata <= 8'h47;
            13'h19F2: rddata <= 8'h38;
            13'h19F3: rddata <= 8'hB7;
            13'h19F4: rddata <= 8'h28;
            13'h19F5: rddata <= 8'h04;
            13'h19F6: rddata <= 8'hAF;
            13'h19F7: rddata <= 8'h32;
            13'h19F8: rddata <= 8'h46;
            13'h19F9: rddata <= 8'h38;
            13'h19FA: rddata <= 8'hC9;
            13'h19FB: rddata <= 8'hD7;
            13'h19FC: rddata <= 8'hE5;
            13'h19FD: rddata <= 8'hCD;
            13'h19FE: rddata <= 8'h18;
            13'h19FF: rddata <= 8'h1A;
            13'h1A00: rddata <= 8'h28;
            13'h1A01: rddata <= 8'h09;
            13'h1A02: rddata <= 8'hF5;
            13'h1A03: rddata <= 8'hCD;
            13'h1A04: rddata <= 8'h4E;
            13'h1A05: rddata <= 8'h0E;
            13'h1A06: rddata <= 8'hF1;
            13'h1A07: rddata <= 8'h5F;
            13'h1A08: rddata <= 8'hCD;
            13'h1A09: rddata <= 8'h19;
            13'h1A0A: rddata <= 8'h10;
            13'h1A0B: rddata <= 8'h21;
            13'h1A0C: rddata <= 8'h6D;
            13'h1A0D: rddata <= 8'h03;
            13'h1A0E: rddata <= 8'h22;
            13'h1A0F: rddata <= 8'hE4;
            13'h1A10: rddata <= 8'h38;
            13'h1A11: rddata <= 8'h3E;
            13'h1A12: rddata <= 8'h01;
            13'h1A13: rddata <= 8'h32;
            13'h1A14: rddata <= 8'hAB;
            13'h1A15: rddata <= 8'h38;
            13'h1A16: rddata <= 8'hE1;
            13'h1A17: rddata <= 8'hC9;
            13'h1A18: rddata <= 8'hE5;
            13'h1A19: rddata <= 8'h21;
            13'h1A1A: rddata <= 8'h0A;
            13'h1A1B: rddata <= 8'h38;
            13'h1A1C: rddata <= 8'h7E;
            13'h1A1D: rddata <= 8'h36;
            13'h1A1E: rddata <= 8'h00;
            13'h1A1F: rddata <= 8'hB7;
            13'h1A20: rddata <= 8'hCC;
            13'h1A21: rddata <= 8'h39;
            13'h1A22: rddata <= 8'h1A;
            13'h1A23: rddata <= 8'hE1;
            13'h1A24: rddata <= 8'hC9;
            13'h1A25: rddata <= 8'hCD;
            13'h1A26: rddata <= 8'h39;
            13'h1A27: rddata <= 8'h1A;
            13'h1A28: rddata <= 8'hC8;
            13'h1A29: rddata <= 8'h32;
            13'h1A2A: rddata <= 8'h0A;
            13'h1A2B: rddata <= 8'h38;
            13'h1A2C: rddata <= 8'hFE;
            13'h1A2D: rddata <= 8'h13;
            13'h1A2E: rddata <= 8'hC0;
            13'h1A2F: rddata <= 8'hAF;
            13'h1A30: rddata <= 8'h32;
            13'h1A31: rddata <= 8'h0A;
            13'h1A32: rddata <= 8'h38;
            13'h1A33: rddata <= 8'hCD;
            13'h1A34: rddata <= 8'h39;
            13'h1A35: rddata <= 8'h1A;
            13'h1A36: rddata <= 8'h28;
            13'h1A37: rddata <= 8'hFB;
            13'h1A38: rddata <= 8'hC9;
            13'h1A39: rddata <= 8'hCD;
            13'h1A3A: rddata <= 8'h7E;
            13'h1A3B: rddata <= 8'h1E;
            13'h1A3C: rddata <= 8'hFE;
            13'h1A3D: rddata <= 8'h03;
            13'h1A3E: rddata <= 8'h20;
            13'h1A3F: rddata <= 8'h0A;
            13'h1A40: rddata <= 8'h3A;
            13'h1A41: rddata <= 8'h5E;
            13'h1A42: rddata <= 8'h38;
            13'h1A43: rddata <= 8'hB7;
            13'h1A44: rddata <= 8'hCC;
            13'h1A45: rddata <= 8'hBE;
            13'h1A46: rddata <= 8'h0B;
            13'h1A47: rddata <= 8'hC3;
            13'h1A48: rddata <= 8'hCE;
            13'h1A49: rddata <= 8'h1F;
            13'h1A4A: rddata <= 8'hB7;
            13'h1A4B: rddata <= 8'hC9;
            13'h1A4C: rddata <= 8'hAF;
            13'h1A4D: rddata <= 8'h18;
            13'h1A4E: rddata <= 8'h02;
            13'h1A4F: rddata <= 8'h3E;
            13'h1A50: rddata <= 8'h01;
            13'h1A51: rddata <= 8'h08;
            13'h1A52: rddata <= 8'hCD;
            13'h1A53: rddata <= 8'h7F;
            13'h1A54: rddata <= 8'h1A;
            13'h1A55: rddata <= 8'hCD;
            13'h1A56: rddata <= 8'h8E;
            13'h1A57: rddata <= 8'h1A;
            13'h1A58: rddata <= 8'h28;
            13'h1A59: rddata <= 8'h02;
            13'h1A5A: rddata <= 8'h36;
            13'h1A5B: rddata <= 8'hA0;
            13'h1A5C: rddata <= 8'h08;
            13'h1A5D: rddata <= 8'hB7;
            13'h1A5E: rddata <= 8'h1A;
            13'h1A5F: rddata <= 8'h20;
            13'h1A60: rddata <= 8'h03;
            13'h1A61: rddata <= 8'h2F;
            13'h1A62: rddata <= 8'hA6;
            13'h1A63: rddata <= 8'h06;
            13'h1A64: rddata <= 8'hB6;
            13'h1A65: rddata <= 8'h77;
            13'h1A66: rddata <= 8'hE1;
            13'h1A67: rddata <= 8'hC9;
            13'h1A68: rddata <= 8'hD7;
            13'h1A69: rddata <= 8'hCD;
            13'h1A6A: rddata <= 8'h7F;
            13'h1A6B: rddata <= 8'h1A;
            13'h1A6C: rddata <= 8'hCD;
            13'h1A6D: rddata <= 8'h8E;
            13'h1A6E: rddata <= 8'h1A;
            13'h1A6F: rddata <= 8'h20;
            13'h1A70: rddata <= 8'h06;
            13'h1A71: rddata <= 8'h1A;
            13'h1A72: rddata <= 8'hA6;
            13'h1A73: rddata <= 8'h16;
            13'h1A74: rddata <= 8'h01;
            13'h1A75: rddata <= 8'h20;
            13'h1A76: rddata <= 8'h02;
            13'h1A77: rddata <= 8'h16;
            13'h1A78: rddata <= 8'h00;
            13'h1A79: rddata <= 8'hAF;
            13'h1A7A: rddata <= 8'hCD;
            13'h1A7B: rddata <= 8'h23;
            13'h1A7C: rddata <= 8'h0B;
            13'h1A7D: rddata <= 8'hE1;
            13'h1A7E: rddata <= 8'hC9;
            13'h1A7F: rddata <= 8'hCF;
            13'h1A80: rddata <= 8'h28;
            13'h1A81: rddata <= 8'hCD;
            13'h1A82: rddata <= 8'hD0;
            13'h1A83: rddata <= 8'h1A;
            13'h1A84: rddata <= 8'hD5;
            13'h1A85: rddata <= 8'hCF;
            13'h1A86: rddata <= 8'h2C;
            13'h1A87: rddata <= 8'hCD;
            13'h1A88: rddata <= 8'hD0;
            13'h1A89: rddata <= 8'h1A;
            13'h1A8A: rddata <= 8'hCF;
            13'h1A8B: rddata <= 8'h29;
            13'h1A8C: rddata <= 8'hC1;
            13'h1A8D: rddata <= 8'hC9;
            13'h1A8E: rddata <= 8'hE3;
            13'h1A8F: rddata <= 8'hE5;
            13'h1A90: rddata <= 8'hC5;
            13'h1A91: rddata <= 8'hD5;
            13'h1A92: rddata <= 8'h21;
            13'h1A93: rddata <= 8'h47;
            13'h1A94: rddata <= 8'h00;
            13'h1A95: rddata <= 8'hE7;
            13'h1A96: rddata <= 8'hDA;
            13'h1A97: rddata <= 8'h97;
            13'h1A98: rddata <= 8'h06;
            13'h1A99: rddata <= 8'h21;
            13'h1A9A: rddata <= 8'h4F;
            13'h1A9B: rddata <= 8'h00;
            13'h1A9C: rddata <= 8'hC5;
            13'h1A9D: rddata <= 8'hD1;
            13'h1A9E: rddata <= 8'hE7;
            13'h1A9F: rddata <= 8'h38;
            13'h1AA0: rddata <= 8'hF5;
            13'h1AA1: rddata <= 8'hD1;
            13'h1AA2: rddata <= 8'hC1;
            13'h1AA3: rddata <= 8'h21;
            13'h1AA4: rddata <= 8'h28;
            13'h1AA5: rddata <= 8'h30;
            13'h1AA6: rddata <= 8'h7B;
            13'h1AA7: rddata <= 8'h11;
            13'h1AA8: rddata <= 8'h28;
            13'h1AA9: rddata <= 8'h00;
            13'h1AAA: rddata <= 8'hFE;
            13'h1AAB: rddata <= 8'h03;
            13'h1AAC: rddata <= 8'h38;
            13'h1AAD: rddata <= 8'h06;
            13'h1AAE: rddata <= 8'h19;
            13'h1AAF: rddata <= 8'h3D;
            13'h1AB0: rddata <= 8'h3D;
            13'h1AB1: rddata <= 8'h3D;
            13'h1AB2: rddata <= 8'h18;
            13'h1AB3: rddata <= 8'hF6;
            13'h1AB4: rddata <= 8'h07;
            13'h1AB5: rddata <= 8'hCB;
            13'h1AB6: rddata <= 8'h29;
            13'h1AB7: rddata <= 8'h30;
            13'h1AB8: rddata <= 8'h01;
            13'h1AB9: rddata <= 8'h3C;
            13'h1ABA: rddata <= 8'h09;
            13'h1ABB: rddata <= 8'h11;
            13'h1ABC: rddata <= 8'hCA;
            13'h1ABD: rddata <= 8'h1A;
            13'h1ABE: rddata <= 8'hB7;
            13'h1ABF: rddata <= 8'h28;
            13'h1AC0: rddata <= 8'h04;
            13'h1AC1: rddata <= 8'h13;
            13'h1AC2: rddata <= 8'h3D;
            13'h1AC3: rddata <= 8'h18;
            13'h1AC4: rddata <= 8'hF9;
            13'h1AC5: rddata <= 8'h7E;
            13'h1AC6: rddata <= 8'hF6;
            13'h1AC7: rddata <= 8'hA0;
            13'h1AC8: rddata <= 8'hAE;
            13'h1AC9: rddata <= 8'hC9;
            13'h1ACA: rddata <= 8'h01;
            13'h1ACB: rddata <= 8'h02;
            13'h1ACC: rddata <= 8'h04;
            13'h1ACD: rddata <= 8'h08;
            13'h1ACE: rddata <= 8'h10;
            13'h1ACF: rddata <= 8'h40;
            13'h1AD0: rddata <= 8'hCD;
            13'h1AD1: rddata <= 8'h85;
            13'h1AD2: rddata <= 8'h09;
            13'h1AD3: rddata <= 8'hC3;
            13'h1AD4: rddata <= 8'h82;
            13'h1AD5: rddata <= 8'h06;
            13'h1AD6: rddata <= 8'hD5;
            13'h1AD7: rddata <= 8'hCD;
            13'h1AD8: rddata <= 8'h7F;
            13'h1AD9: rddata <= 8'h1A;
            13'h1ADA: rddata <= 8'hE5;
            13'h1ADB: rddata <= 8'hCD;
            13'h1ADC: rddata <= 8'h64;
            13'h1ADD: rddata <= 8'h1E;
            13'h1ADE: rddata <= 8'hE1;
            13'h1ADF: rddata <= 8'hD1;
            13'h1AE0: rddata <= 8'hC9;
            13'h1AE1: rddata <= 8'h3E;
            13'h1AE2: rddata <= 8'h0D;
            13'h1AE3: rddata <= 8'hCD;
            13'h1AE4: rddata <= 8'hE8;
            13'h1AE5: rddata <= 8'h1A;
            13'h1AE6: rddata <= 8'h3E;
            13'h1AE7: rddata <= 8'h0A;
            13'h1AE8: rddata <= 8'hF7;
            13'h1AE9: rddata <= 8'h11;
            13'h1AEA: rddata <= 8'hF5;
            13'h1AEB: rddata <= 8'hF5;
            13'h1AEC: rddata <= 8'hD9;
            13'h1AED: rddata <= 8'hDB;
            13'h1AEE: rddata <= 8'hFE;
            13'h1AEF: rddata <= 8'hE6;
            13'h1AF0: rddata <= 8'h01;
            13'h1AF1: rddata <= 8'h28;
            13'h1AF2: rddata <= 8'hFA;
            13'h1AF3: rddata <= 8'hCD;
            13'h1AF4: rddata <= 8'h08;
            13'h1AF5: rddata <= 8'h1B;
            13'h1AF6: rddata <= 8'h1E;
            13'h1AF7: rddata <= 8'h08;
            13'h1AF8: rddata <= 8'hF1;
            13'h1AF9: rddata <= 8'hCD;
            13'h1AFA: rddata <= 8'h0A;
            13'h1AFB: rddata <= 8'h1B;
            13'h1AFC: rddata <= 8'h0F;
            13'h1AFD: rddata <= 8'h1D;
            13'h1AFE: rddata <= 8'h20;
            13'h1AFF: rddata <= 8'hF9;
            13'h1B00: rddata <= 8'h3E;
            13'h1B01: rddata <= 8'h01;
            13'h1B02: rddata <= 8'hCD;
            13'h1B03: rddata <= 8'h0A;
            13'h1B04: rddata <= 8'h1B;
            13'h1B05: rddata <= 8'hD9;
            13'h1B06: rddata <= 8'hF1;
            13'h1B07: rddata <= 8'hC9;
            13'h1B08: rddata <= 8'h3E;
            13'h1B09: rddata <= 8'h00;
            13'h1B0A: rddata <= 8'hD3;
            13'h1B0B: rddata <= 8'hFE;
            13'h1B0C: rddata <= 8'h26;
            13'h1B0D: rddata <= 8'hB1;
            13'h1B0E: rddata <= 8'h25;
            13'h1B0F: rddata <= 8'h20;
            13'h1B10: rddata <= 8'hFD;
            13'h1B11: rddata <= 8'h00;
            13'h1B12: rddata <= 8'h00;
            13'h1B13: rddata <= 8'h00;
            13'h1B14: rddata <= 8'hC9;
            13'h1B15: rddata <= 8'hE5;
            13'h1B16: rddata <= 8'hD5;
            13'h1B17: rddata <= 8'hCD;
            13'h1B18: rddata <= 8'hE1;
            13'h1B19: rddata <= 8'h1A;
            13'h1B1A: rddata <= 8'h21;
            13'h1B1B: rddata <= 8'h28;
            13'h1B1C: rddata <= 8'h30;
            13'h1B1D: rddata <= 8'h11;
            13'h1B1E: rddata <= 8'hE8;
            13'h1B1F: rddata <= 8'h33;
            13'h1B20: rddata <= 8'h7E;
            13'h1B21: rddata <= 8'hCD;
            13'h1B22: rddata <= 8'hE8;
            13'h1B23: rddata <= 8'h1A;
            13'h1B24: rddata <= 8'h23;
            13'h1B25: rddata <= 8'hE7;
            13'h1B26: rddata <= 8'h38;
            13'h1B27: rddata <= 8'hF8;
            13'h1B28: rddata <= 8'hCD;
            13'h1B29: rddata <= 8'hE1;
            13'h1B2A: rddata <= 8'h1A;
            13'h1B2B: rddata <= 8'hD1;
            13'h1B2C: rddata <= 8'hE1;
            13'h1B2D: rddata <= 8'hC9;
            13'h1B2E: rddata <= 8'hE5;
            13'h1B2F: rddata <= 8'hD5;
            13'h1B30: rddata <= 8'hC5;
            13'h1B31: rddata <= 8'h21;
            13'h1B32: rddata <= 8'hE8;
            13'h1B33: rddata <= 8'h1B;
            13'h1B34: rddata <= 8'hF5;
            13'h1B35: rddata <= 8'hCD;
            13'h1B36: rddata <= 8'h9D;
            13'h1B37: rddata <= 8'h0E;
            13'h1B38: rddata <= 8'h21;
            13'h1B39: rddata <= 8'hB5;
            13'h1B3A: rddata <= 8'h00;
            13'h1B3B: rddata <= 8'hCD;
            13'h1B3C: rddata <= 8'h9D;
            13'h1B3D: rddata <= 8'h0E;
            13'h1B3E: rddata <= 8'hCD;
            13'h1B3F: rddata <= 8'h7E;
            13'h1B40: rddata <= 8'h1E;
            13'h1B41: rddata <= 8'hFE;
            13'h1B42: rddata <= 8'h0D;
            13'h1B43: rddata <= 8'h20;
            13'h1B44: rddata <= 8'hF9;
            13'h1B45: rddata <= 8'hCD;
            13'h1B46: rddata <= 8'hEA;
            13'h1B47: rddata <= 8'h19;
            13'h1B48: rddata <= 8'hF1;
            13'h1B49: rddata <= 8'hC1;
            13'h1B4A: rddata <= 8'hD1;
            13'h1B4B: rddata <= 8'hE1;
            13'h1B4C: rddata <= 8'hC9;
            13'h1B4D: rddata <= 8'hD9;
            13'h1B4E: rddata <= 8'h0E;
            13'h1B4F: rddata <= 8'hFC;
            13'h1B50: rddata <= 8'hCD;
            13'h1B51: rddata <= 8'h62;
            13'h1B52: rddata <= 8'h1B;
            13'h1B53: rddata <= 8'h38;
            13'h1B54: rddata <= 8'hFB;
            13'h1B55: rddata <= 8'h26;
            13'h1B56: rddata <= 8'h08;
            13'h1B57: rddata <= 8'hCD;
            13'h1B58: rddata <= 8'h62;
            13'h1B59: rddata <= 8'h1B;
            13'h1B5A: rddata <= 8'hCB;
            13'h1B5B: rddata <= 8'h15;
            13'h1B5C: rddata <= 8'h25;
            13'h1B5D: rddata <= 8'h20;
            13'h1B5E: rddata <= 8'hF8;
            13'h1B5F: rddata <= 8'h7D;
            13'h1B60: rddata <= 8'hD9;
            13'h1B61: rddata <= 8'hC9;
            13'h1B62: rddata <= 8'hED;
            13'h1B63: rddata <= 8'h78;
            13'h1B64: rddata <= 8'h1F;
            13'h1B65: rddata <= 8'h38;
            13'h1B66: rddata <= 8'hFB;
            13'h1B67: rddata <= 8'hED;
            13'h1B68: rddata <= 8'h78;
            13'h1B69: rddata <= 8'h1F;
            13'h1B6A: rddata <= 8'h30;
            13'h1B6B: rddata <= 8'hFB;
            13'h1B6C: rddata <= 8'hAF;
            13'h1B6D: rddata <= 8'h3C;
            13'h1B6E: rddata <= 8'hED;
            13'h1B6F: rddata <= 8'h40;
            13'h1B70: rddata <= 8'hCB;
            13'h1B71: rddata <= 8'h18;
            13'h1B72: rddata <= 8'h38;
            13'h1B73: rddata <= 8'hF9;
            13'h1B74: rddata <= 8'h3C;
            13'h1B75: rddata <= 8'hED;
            13'h1B76: rddata <= 8'h40;
            13'h1B77: rddata <= 8'hCB;
            13'h1B78: rddata <= 8'h18;
            13'h1B79: rddata <= 8'h30;
            13'h1B7A: rddata <= 8'hF9;
            13'h1B7B: rddata <= 8'hFE;
            13'h1B7C: rddata <= 8'h49;
            13'h1B7D: rddata <= 8'hC9;
            13'h1B7E: rddata <= 8'hC9;
            13'h1B7F: rddata <= 8'hE5;
            13'h1B80: rddata <= 8'hD5;
            13'h1B81: rddata <= 8'hC5;
            13'h1B82: rddata <= 8'h21;
            13'h1B83: rddata <= 8'hF7;
            13'h1B84: rddata <= 8'h1B;
            13'h1B85: rddata <= 8'h18;
            13'h1B86: rddata <= 8'hAD;
            13'h1B87: rddata <= 8'hCD;
            13'h1B88: rddata <= 8'h8A;
            13'h1B89: rddata <= 8'h1B;
            13'h1B8A: rddata <= 8'hF5;
            13'h1B8B: rddata <= 8'hD9;
            13'h1B8C: rddata <= 8'h0E;
            13'h1B8D: rddata <= 8'hFC;
            13'h1B8E: rddata <= 8'hF5;
            13'h1B8F: rddata <= 8'hAF;
            13'h1B90: rddata <= 8'h1E;
            13'h1B91: rddata <= 8'h01;
            13'h1B92: rddata <= 8'hCD;
            13'h1B93: rddata <= 8'hA5;
            13'h1B94: rddata <= 8'h1B;
            13'h1B95: rddata <= 8'hF1;
            13'h1B96: rddata <= 8'h1E;
            13'h1B97: rddata <= 8'h08;
            13'h1B98: rddata <= 8'hCD;
            13'h1B99: rddata <= 8'hA5;
            13'h1B9A: rddata <= 8'h1B;
            13'h1B9B: rddata <= 8'h3E;
            13'h1B9C: rddata <= 8'hFF;
            13'h1B9D: rddata <= 8'h1E;
            13'h1B9E: rddata <= 8'h02;
            13'h1B9F: rddata <= 8'hCD;
            13'h1BA0: rddata <= 8'hA5;
            13'h1BA1: rddata <= 8'h1B;
            13'h1BA2: rddata <= 8'hD9;
            13'h1BA3: rddata <= 8'hF1;
            13'h1BA4: rddata <= 8'hC9;
            13'h1BA5: rddata <= 8'h17;
            13'h1BA6: rddata <= 8'h2E;
            13'h1BA7: rddata <= 8'h40;
            13'h1BA8: rddata <= 8'h38;
            13'h1BA9: rddata <= 8'h02;
            13'h1BAA: rddata <= 8'h2E;
            13'h1BAB: rddata <= 8'h80;
            13'h1BAC: rddata <= 8'h06;
            13'h1BAD: rddata <= 8'h04;
            13'h1BAE: rddata <= 8'hED;
            13'h1BAF: rddata <= 8'h41;
            13'h1BB0: rddata <= 8'h65;
            13'h1BB1: rddata <= 8'h25;
            13'h1BB2: rddata <= 8'h20;
            13'h1BB3: rddata <= 8'hFD;
            13'h1BB4: rddata <= 8'h05;
            13'h1BB5: rddata <= 8'h20;
            13'h1BB6: rddata <= 8'hF7;
            13'h1BB7: rddata <= 8'h1D;
            13'h1BB8: rddata <= 8'h20;
            13'h1BB9: rddata <= 8'hEB;
            13'h1BBA: rddata <= 8'hC9;
            13'h1BBB: rddata <= 8'hC9;
            13'h1BBC: rddata <= 8'hF5;
            13'h1BBD: rddata <= 8'hC5;
            13'h1BBE: rddata <= 8'h06;
            13'h1BBF: rddata <= 8'h0C;
            13'h1BC0: rddata <= 8'h3E;
            13'h1BC1: rddata <= 8'hFF;
            13'h1BC2: rddata <= 8'hCD;
            13'h1BC3: rddata <= 8'h8A;
            13'h1BC4: rddata <= 8'h1B;
            13'h1BC5: rddata <= 8'h10;
            13'h1BC6: rddata <= 8'hF9;
            13'h1BC7: rddata <= 8'hAF;
            13'h1BC8: rddata <= 8'hCD;
            13'h1BC9: rddata <= 8'h8A;
            13'h1BCA: rddata <= 8'h1B;
            13'h1BCB: rddata <= 8'hC1;
            13'h1BCC: rddata <= 8'hF1;
            13'h1BCD: rddata <= 8'hC9;
            13'h1BCE: rddata <= 8'hF5;
            13'h1BCF: rddata <= 8'hC5;
            13'h1BD0: rddata <= 8'h06;
            13'h1BD1: rddata <= 8'h06;
            13'h1BD2: rddata <= 8'hCD;
            13'h1BD3: rddata <= 8'h4D;
            13'h1BD4: rddata <= 8'h1B;
            13'h1BD5: rddata <= 8'h3C;
            13'h1BD6: rddata <= 8'h20;
            13'h1BD7: rddata <= 8'hF8;
            13'h1BD8: rddata <= 8'h10;
            13'h1BD9: rddata <= 8'hF8;
            13'h1BDA: rddata <= 8'hCD;
            13'h1BDB: rddata <= 8'h4D;
            13'h1BDC: rddata <= 8'h1B;
            13'h1BDD: rddata <= 8'hB7;
            13'h1BDE: rddata <= 8'h28;
            13'h1BDF: rddata <= 8'h05;
            13'h1BE0: rddata <= 8'h3C;
            13'h1BE1: rddata <= 8'h28;
            13'h1BE2: rddata <= 8'hF7;
            13'h1BE3: rddata <= 8'h18;
            13'h1BE4: rddata <= 8'hEB;
            13'h1BE5: rddata <= 8'hC1;
            13'h1BE6: rddata <= 8'hF1;
            13'h1BE7: rddata <= 8'hC9;
            13'h1BE8: rddata <= 8'h50;
            13'h1BE9: rddata <= 8'h72;
            13'h1BEA: rddata <= 8'h65;
            13'h1BEB: rddata <= 8'h73;
            13'h1BEC: rddata <= 8'h73;
            13'h1BED: rddata <= 8'h20;
            13'h1BEE: rddata <= 8'h3C;
            13'h1BEF: rddata <= 8'h50;
            13'h1BF0: rddata <= 8'h4C;
            13'h1BF1: rddata <= 8'h41;
            13'h1BF2: rddata <= 8'h59;
            13'h1BF3: rddata <= 8'h3E;
            13'h1BF4: rddata <= 8'h0D;
            13'h1BF5: rddata <= 8'h0A;
            13'h1BF6: rddata <= 8'h00;
            13'h1BF7: rddata <= 8'h50;
            13'h1BF8: rddata <= 8'h72;
            13'h1BF9: rddata <= 8'h65;
            13'h1BFA: rddata <= 8'h73;
            13'h1BFB: rddata <= 8'h73;
            13'h1BFC: rddata <= 8'h20;
            13'h1BFD: rddata <= 8'h3C;
            13'h1BFE: rddata <= 8'h52;
            13'h1BFF: rddata <= 8'h45;
            13'h1C00: rddata <= 8'h43;
            13'h1C01: rddata <= 8'h4F;
            13'h1C02: rddata <= 8'h52;
            13'h1C03: rddata <= 8'h44;
            13'h1C04: rddata <= 8'h3E;
            13'h1C05: rddata <= 8'h0D;
            13'h1C06: rddata <= 8'h0A;
            13'h1C07: rddata <= 8'h00;
            13'h1C08: rddata <= 8'hF7;
            13'h1C09: rddata <= 8'h15;
            13'h1C0A: rddata <= 8'hFE;
            13'h1C0B: rddata <= 8'hAA;
            13'h1C0C: rddata <= 8'hCA;
            13'h1C0D: rddata <= 8'h62;
            13'h1C0E: rddata <= 8'h0C;
            13'h1C0F: rddata <= 8'hCD;
            13'h1C10: rddata <= 8'hB8;
            13'h1C11: rddata <= 8'h1C;
            13'h1C12: rddata <= 8'hE5;
            13'h1C13: rddata <= 8'hCD;
            13'h1C14: rddata <= 8'h25;
            13'h1C15: rddata <= 8'h1D;
            13'h1C16: rddata <= 8'h2A;
            13'h1C17: rddata <= 8'h4F;
            13'h1C18: rddata <= 8'h38;
            13'h1C19: rddata <= 8'hCD;
            13'h1C1A: rddata <= 8'h38;
            13'h1C1B: rddata <= 8'h1D;
            13'h1C1C: rddata <= 8'h06;
            13'h1C1D: rddata <= 8'h0F;
            13'h1C1E: rddata <= 8'hAF;
            13'h1C1F: rddata <= 8'hCD;
            13'h1C20: rddata <= 8'h8A;
            13'h1C21: rddata <= 8'h1B;
            13'h1C22: rddata <= 8'h10;
            13'h1C23: rddata <= 8'hFB;
            13'h1C24: rddata <= 8'h01;
            13'h1C25: rddata <= 8'h40;
            13'h1C26: rddata <= 8'h1F;
            13'h1C27: rddata <= 8'hCD;
            13'h1C28: rddata <= 8'h4B;
            13'h1C29: rddata <= 8'h1D;
            13'h1C2A: rddata <= 8'hE1;
            13'h1C2B: rddata <= 8'hC9;
            13'h1C2C: rddata <= 8'hF7;
            13'h1C2D: rddata <= 8'h14;
            13'h1C2E: rddata <= 8'hFE;
            13'h1C2F: rddata <= 8'hAA;
            13'h1C30: rddata <= 8'hCA;
            13'h1C31: rddata <= 8'h63;
            13'h1C32: rddata <= 8'h0C;
            13'h1C33: rddata <= 8'hD6;
            13'h1C34: rddata <= 8'h95;
            13'h1C35: rddata <= 8'h28;
            13'h1C36: rddata <= 8'h02;
            13'h1C37: rddata <= 8'hAF;
            13'h1C38: rddata <= 8'h01;
            13'h1C39: rddata <= 8'h2F;
            13'h1C3A: rddata <= 8'h23;
            13'h1C3B: rddata <= 8'hFE;
            13'h1C3C: rddata <= 8'h01;
            13'h1C3D: rddata <= 8'hF5;
            13'h1C3E: rddata <= 8'h3E;
            13'h1C3F: rddata <= 8'hFF;
            13'h1C40: rddata <= 8'h32;
            13'h1C41: rddata <= 8'h5E;
            13'h1C42: rddata <= 8'h38;
            13'h1C43: rddata <= 8'hCD;
            13'h1C44: rddata <= 8'hB1;
            13'h1C45: rddata <= 8'h1C;
            13'h1C46: rddata <= 8'hAF;
            13'h1C47: rddata <= 8'h32;
            13'h1C48: rddata <= 8'h5D;
            13'h1C49: rddata <= 8'h38;
            13'h1C4A: rddata <= 8'hD5;
            13'h1C4B: rddata <= 8'hCD;
            13'h1C4C: rddata <= 8'h2E;
            13'h1C4D: rddata <= 8'h1B;
            13'h1C4E: rddata <= 8'hCD;
            13'h1C4F: rddata <= 8'hD9;
            13'h1C50: rddata <= 8'h1C;
            13'h1C51: rddata <= 8'h21;
            13'h1C52: rddata <= 8'h57;
            13'h1C53: rddata <= 8'h38;
            13'h1C54: rddata <= 8'hCD;
            13'h1C55: rddata <= 8'hED;
            13'h1C56: rddata <= 8'h1C;
            13'h1C57: rddata <= 8'hD1;
            13'h1C58: rddata <= 8'h28;
            13'h1C59: rddata <= 8'h12;
            13'h1C5A: rddata <= 8'h21;
            13'h1C5B: rddata <= 8'h06;
            13'h1C5C: rddata <= 8'h1D;
            13'h1C5D: rddata <= 8'hCD;
            13'h1C5E: rddata <= 8'h0D;
            13'h1C5F: rddata <= 8'h1D;
            13'h1C60: rddata <= 8'h06;
            13'h1C61: rddata <= 8'h0A;
            13'h1C62: rddata <= 8'hCD;
            13'h1C63: rddata <= 8'h4D;
            13'h1C64: rddata <= 8'h1B;
            13'h1C65: rddata <= 8'hB7;
            13'h1C66: rddata <= 8'h20;
            13'h1C67: rddata <= 8'hF8;
            13'h1C68: rddata <= 8'h10;
            13'h1C69: rddata <= 8'hF8;
            13'h1C6A: rddata <= 8'h18;
            13'h1C6B: rddata <= 8'hDA;
            13'h1C6C: rddata <= 8'h21;
            13'h1C6D: rddata <= 8'hFE;
            13'h1C6E: rddata <= 8'h1C;
            13'h1C6F: rddata <= 8'hCD;
            13'h1C70: rddata <= 8'h0D;
            13'h1C71: rddata <= 8'h1D;
            13'h1C72: rddata <= 8'hF1;
            13'h1C73: rddata <= 8'h32;
            13'h1C74: rddata <= 8'hE4;
            13'h1C75: rddata <= 8'h38;
            13'h1C76: rddata <= 8'hDC;
            13'h1C77: rddata <= 8'hBE;
            13'h1C78: rddata <= 8'h0B;
            13'h1C79: rddata <= 8'h3A;
            13'h1C7A: rddata <= 8'hE4;
            13'h1C7B: rddata <= 8'h38;
            13'h1C7C: rddata <= 8'hFE;
            13'h1C7D: rddata <= 8'h01;
            13'h1C7E: rddata <= 8'h32;
            13'h1C7F: rddata <= 8'h5E;
            13'h1C80: rddata <= 8'h38;
            13'h1C81: rddata <= 8'h2A;
            13'h1C82: rddata <= 8'h4F;
            13'h1C83: rddata <= 8'h38;
            13'h1C84: rddata <= 8'hCD;
            13'h1C85: rddata <= 8'h51;
            13'h1C86: rddata <= 8'h1D;
            13'h1C87: rddata <= 8'h20;
            13'h1C88: rddata <= 8'h11;
            13'h1C89: rddata <= 8'h22;
            13'h1C8A: rddata <= 8'hD6;
            13'h1C8B: rddata <= 8'h38;
            13'h1C8C: rddata <= 8'h21;
            13'h1C8D: rddata <= 8'h6E;
            13'h1C8E: rddata <= 8'h03;
            13'h1C8F: rddata <= 8'hCD;
            13'h1C90: rddata <= 8'h9D;
            13'h1C91: rddata <= 8'h0E;
            13'h1C92: rddata <= 8'h3E;
            13'h1C93: rddata <= 8'hFF;
            13'h1C94: rddata <= 8'h32;
            13'h1C95: rddata <= 8'h5E;
            13'h1C96: rddata <= 8'h38;
            13'h1C97: rddata <= 8'hC3;
            13'h1C98: rddata <= 8'h80;
            13'h1C99: rddata <= 8'h04;
            13'h1C9A: rddata <= 8'h23;
            13'h1C9B: rddata <= 8'hEB;
            13'h1C9C: rddata <= 8'h2A;
            13'h1C9D: rddata <= 8'hD6;
            13'h1C9E: rddata <= 8'h38;
            13'h1C9F: rddata <= 8'hE7;
            13'h1CA0: rddata <= 8'h38;
            13'h1CA1: rddata <= 8'hEA;
            13'h1CA2: rddata <= 8'h21;
            13'h1CA3: rddata <= 8'hAB;
            13'h1CA4: rddata <= 8'h1C;
            13'h1CA5: rddata <= 8'hCD;
            13'h1CA6: rddata <= 8'h9D;
            13'h1CA7: rddata <= 8'h0E;
            13'h1CA8: rddata <= 8'hC3;
            13'h1CA9: rddata <= 8'h01;
            13'h1CAA: rddata <= 8'h04;
            13'h1CAB: rddata <= 8'h42;
            13'h1CAC: rddata <= 8'h61;
            13'h1CAD: rddata <= 8'h64;
            13'h1CAE: rddata <= 8'h0D;
            13'h1CAF: rddata <= 8'h0A;
            13'h1CB0: rddata <= 8'h00;
            13'h1CB1: rddata <= 8'hAF;
            13'h1CB2: rddata <= 8'h32;
            13'h1CB3: rddata <= 8'h51;
            13'h1CB4: rddata <= 8'h38;
            13'h1CB5: rddata <= 8'h2B;
            13'h1CB6: rddata <= 8'hD7;
            13'h1CB7: rddata <= 8'hC8;
            13'h1CB8: rddata <= 8'hCD;
            13'h1CB9: rddata <= 8'h85;
            13'h1CBA: rddata <= 8'h09;
            13'h1CBB: rddata <= 8'hE5;
            13'h1CBC: rddata <= 8'hCD;
            13'h1CBD: rddata <= 8'h06;
            13'h1CBE: rddata <= 8'h10;
            13'h1CBF: rddata <= 8'h2B;
            13'h1CC0: rddata <= 8'h2B;
            13'h1CC1: rddata <= 8'h2B;
            13'h1CC2: rddata <= 8'h46;
            13'h1CC3: rddata <= 8'h0E;
            13'h1CC4: rddata <= 8'h06;
            13'h1CC5: rddata <= 8'h21;
            13'h1CC6: rddata <= 8'h51;
            13'h1CC7: rddata <= 8'h38;
            13'h1CC8: rddata <= 8'h1A;
            13'h1CC9: rddata <= 8'h77;
            13'h1CCA: rddata <= 8'h23;
            13'h1CCB: rddata <= 8'h13;
            13'h1CCC: rddata <= 8'h0D;
            13'h1CCD: rddata <= 8'h28;
            13'h1CCE: rddata <= 8'h08;
            13'h1CCF: rddata <= 8'h10;
            13'h1CD0: rddata <= 8'hF7;
            13'h1CD1: rddata <= 8'h41;
            13'h1CD2: rddata <= 8'h36;
            13'h1CD3: rddata <= 8'h00;
            13'h1CD4: rddata <= 8'h23;
            13'h1CD5: rddata <= 8'h10;
            13'h1CD6: rddata <= 8'hFB;
            13'h1CD7: rddata <= 8'hE1;
            13'h1CD8: rddata <= 8'hC9;
            13'h1CD9: rddata <= 8'hCD;
            13'h1CDA: rddata <= 8'hCE;
            13'h1CDB: rddata <= 8'h1B;
            13'h1CDC: rddata <= 8'hAF;
            13'h1CDD: rddata <= 8'h32;
            13'h1CDE: rddata <= 8'h5D;
            13'h1CDF: rddata <= 8'h38;
            13'h1CE0: rddata <= 8'h21;
            13'h1CE1: rddata <= 8'h57;
            13'h1CE2: rddata <= 8'h38;
            13'h1CE3: rddata <= 8'h06;
            13'h1CE4: rddata <= 8'h06;
            13'h1CE5: rddata <= 8'hCD;
            13'h1CE6: rddata <= 8'h4D;
            13'h1CE7: rddata <= 8'h1B;
            13'h1CE8: rddata <= 8'h77;
            13'h1CE9: rddata <= 8'h23;
            13'h1CEA: rddata <= 8'h10;
            13'h1CEB: rddata <= 8'hF9;
            13'h1CEC: rddata <= 8'hC9;
            13'h1CED: rddata <= 8'h01;
            13'h1CEE: rddata <= 8'h51;
            13'h1CEF: rddata <= 8'h38;
            13'h1CF0: rddata <= 8'h1E;
            13'h1CF1: rddata <= 8'h06;
            13'h1CF2: rddata <= 8'h0A;
            13'h1CF3: rddata <= 8'hB7;
            13'h1CF4: rddata <= 8'hC8;
            13'h1CF5: rddata <= 8'h0A;
            13'h1CF6: rddata <= 8'hBE;
            13'h1CF7: rddata <= 8'h23;
            13'h1CF8: rddata <= 8'h03;
            13'h1CF9: rddata <= 8'hC0;
            13'h1CFA: rddata <= 8'h1D;
            13'h1CFB: rddata <= 8'h20;
            13'h1CFC: rddata <= 8'hF8;
            13'h1CFD: rddata <= 8'hC9;
            13'h1CFE: rddata <= 8'h46;
            13'h1CFF: rddata <= 8'h6F;
            13'h1D00: rddata <= 8'h75;
            13'h1D01: rddata <= 8'h6E;
            13'h1D02: rddata <= 8'h64;
            13'h1D03: rddata <= 8'h3A;
            13'h1D04: rddata <= 8'h20;
            13'h1D05: rddata <= 8'h00;
            13'h1D06: rddata <= 8'h53;
            13'h1D07: rddata <= 8'h6B;
            13'h1D08: rddata <= 8'h69;
            13'h1D09: rddata <= 8'h70;
            13'h1D0A: rddata <= 8'h3A;
            13'h1D0B: rddata <= 8'h20;
            13'h1D0C: rddata <= 8'h00;
            13'h1D0D: rddata <= 8'hD5;
            13'h1D0E: rddata <= 8'hF5;
            13'h1D0F: rddata <= 8'hCD;
            13'h1D10: rddata <= 8'h9D;
            13'h1D11: rddata <= 8'h0E;
            13'h1D12: rddata <= 8'h21;
            13'h1D13: rddata <= 8'h57;
            13'h1D14: rddata <= 8'h38;
            13'h1D15: rddata <= 8'h06;
            13'h1D16: rddata <= 8'h06;
            13'h1D17: rddata <= 8'h7E;
            13'h1D18: rddata <= 8'h23;
            13'h1D19: rddata <= 8'hB7;
            13'h1D1A: rddata <= 8'h28;
            13'h1D1B: rddata <= 8'h01;
            13'h1D1C: rddata <= 8'hDF;
            13'h1D1D: rddata <= 8'h10;
            13'h1D1E: rddata <= 8'hF8;
            13'h1D1F: rddata <= 8'hCD;
            13'h1D20: rddata <= 8'hEA;
            13'h1D21: rddata <= 8'h19;
            13'h1D22: rddata <= 8'hF1;
            13'h1D23: rddata <= 8'hD1;
            13'h1D24: rddata <= 8'hC9;
            13'h1D25: rddata <= 8'hCD;
            13'h1D26: rddata <= 8'h7F;
            13'h1D27: rddata <= 8'h1B;
            13'h1D28: rddata <= 8'hCD;
            13'h1D29: rddata <= 8'hBC;
            13'h1D2A: rddata <= 8'h1B;
            13'h1D2B: rddata <= 8'h06;
            13'h1D2C: rddata <= 8'h06;
            13'h1D2D: rddata <= 8'h21;
            13'h1D2E: rddata <= 8'h51;
            13'h1D2F: rddata <= 8'h38;
            13'h1D30: rddata <= 8'h7E;
            13'h1D31: rddata <= 8'h23;
            13'h1D32: rddata <= 8'hCD;
            13'h1D33: rddata <= 8'h8A;
            13'h1D34: rddata <= 8'h1B;
            13'h1D35: rddata <= 8'h10;
            13'h1D36: rddata <= 8'hF9;
            13'h1D37: rddata <= 8'hC9;
            13'h1D38: rddata <= 8'hCD;
            13'h1D39: rddata <= 8'hBC;
            13'h1D3A: rddata <= 8'h1B;
            13'h1D3B: rddata <= 8'hEB;
            13'h1D3C: rddata <= 8'h2A;
            13'h1D3D: rddata <= 8'hD6;
            13'h1D3E: rddata <= 8'h38;
            13'h1D3F: rddata <= 8'h1A;
            13'h1D40: rddata <= 8'h13;
            13'h1D41: rddata <= 8'hCD;
            13'h1D42: rddata <= 8'h8A;
            13'h1D43: rddata <= 8'h1B;
            13'h1D44: rddata <= 8'hE7;
            13'h1D45: rddata <= 8'h20;
            13'h1D46: rddata <= 8'hF8;
            13'h1D47: rddata <= 8'hC9;
            13'h1D48: rddata <= 8'h01;
            13'h1D49: rddata <= 8'h00;
            13'h1D4A: rddata <= 8'h00;
            13'h1D4B: rddata <= 8'h0B;
            13'h1D4C: rddata <= 8'h78;
            13'h1D4D: rddata <= 8'hB1;
            13'h1D4E: rddata <= 8'h20;
            13'h1D4F: rddata <= 8'hFB;
            13'h1D50: rddata <= 8'hC9;
            13'h1D51: rddata <= 8'hCD;
            13'h1D52: rddata <= 8'hCE;
            13'h1D53: rddata <= 8'h1B;
            13'h1D54: rddata <= 8'h3E;
            13'h1D55: rddata <= 8'hFF;
            13'h1D56: rddata <= 8'h32;
            13'h1D57: rddata <= 8'h5D;
            13'h1D58: rddata <= 8'h38;
            13'h1D59: rddata <= 8'h9F;
            13'h1D5A: rddata <= 8'h2F;
            13'h1D5B: rddata <= 8'h57;
            13'h1D5C: rddata <= 8'h06;
            13'h1D5D: rddata <= 8'h0A;
            13'h1D5E: rddata <= 8'hCD;
            13'h1D5F: rddata <= 8'h4D;
            13'h1D60: rddata <= 8'h1B;
            13'h1D61: rddata <= 8'h5F;
            13'h1D62: rddata <= 8'h96;
            13'h1D63: rddata <= 8'hA2;
            13'h1D64: rddata <= 8'hC0;
            13'h1D65: rddata <= 8'h73;
            13'h1D66: rddata <= 8'hCD;
            13'h1D67: rddata <= 8'hA9;
            13'h1D68: rddata <= 8'h0B;
            13'h1D69: rddata <= 8'h7E;
            13'h1D6A: rddata <= 8'hB7;
            13'h1D6B: rddata <= 8'h23;
            13'h1D6C: rddata <= 8'h20;
            13'h1D6D: rddata <= 8'hEE;
            13'h1D6E: rddata <= 8'h10;
            13'h1D6F: rddata <= 8'hEE;
            13'h1D70: rddata <= 8'hAF;
            13'h1D71: rddata <= 8'hC9;
            13'h1D72: rddata <= 8'hF7;
            13'h1D73: rddata <= 8'h13;
            13'h1D74: rddata <= 8'hF5;
            13'h1D75: rddata <= 8'hFE;
            13'h1D76: rddata <= 8'h0A;
            13'h1D77: rddata <= 8'h28;
            13'h1D78: rddata <= 8'h1A;
            13'h1D79: rddata <= 8'h3A;
            13'h1D7A: rddata <= 8'h00;
            13'h1D7B: rddata <= 8'h38;
            13'h1D7C: rddata <= 8'hB7;
            13'h1D7D: rddata <= 8'h20;
            13'h1D7E: rddata <= 8'h14;
            13'h1D7F: rddata <= 8'h3A;
            13'h1D80: rddata <= 8'h08;
            13'h1D81: rddata <= 8'h38;
            13'h1D82: rddata <= 8'hB7;
            13'h1D83: rddata <= 8'h28;
            13'h1D84: rddata <= 8'h0E;
            13'h1D85: rddata <= 8'h3D;
            13'h1D86: rddata <= 8'h32;
            13'h1D87: rddata <= 8'h08;
            13'h1D88: rddata <= 8'h38;
            13'h1D89: rddata <= 8'h20;
            13'h1D8A: rddata <= 8'h08;
            13'h1D8B: rddata <= 8'h3E;
            13'h1D8C: rddata <= 8'h17;
            13'h1D8D: rddata <= 8'h32;
            13'h1D8E: rddata <= 8'h08;
            13'h1D8F: rddata <= 8'h38;
            13'h1D90: rddata <= 8'hCD;
            13'h1D91: rddata <= 8'h2F;
            13'h1D92: rddata <= 8'h1A;
            13'h1D93: rddata <= 8'hF1;
            13'h1D94: rddata <= 8'hF5;
            13'h1D95: rddata <= 8'hD9;
            13'h1D96: rddata <= 8'hFE;
            13'h1D97: rddata <= 8'h07;
            13'h1D98: rddata <= 8'hCA;
            13'h1D99: rddata <= 8'h14;
            13'h1D9A: rddata <= 8'h1E;
            13'h1D9B: rddata <= 8'hFE;
            13'h1D9C: rddata <= 8'h0B;
            13'h1D9D: rddata <= 8'hCA;
            13'h1D9E: rddata <= 8'h45;
            13'h1D9F: rddata <= 8'h1E;
            13'h1DA0: rddata <= 8'h5F;
            13'h1DA1: rddata <= 8'h2A;
            13'h1DA2: rddata <= 8'h01;
            13'h1DA3: rddata <= 8'h38;
            13'h1DA4: rddata <= 8'h3A;
            13'h1DA5: rddata <= 8'h0D;
            13'h1DA6: rddata <= 8'h38;
            13'h1DA7: rddata <= 8'h77;
            13'h1DA8: rddata <= 8'h7B;
            13'h1DA9: rddata <= 8'hFE;
            13'h1DAA: rddata <= 8'h08;
            13'h1DAB: rddata <= 8'h28;
            13'h1DAC: rddata <= 8'h30;
            13'h1DAD: rddata <= 8'hFE;
            13'h1DAE: rddata <= 8'h0D;
            13'h1DAF: rddata <= 8'h28;
            13'h1DB0: rddata <= 8'h0D;
            13'h1DB1: rddata <= 8'hFE;
            13'h1DB2: rddata <= 8'h0A;
            13'h1DB3: rddata <= 8'h28;
            13'h1DB4: rddata <= 8'h13;
            13'h1DB5: rddata <= 8'h2A;
            13'h1DB6: rddata <= 8'h01;
            13'h1DB7: rddata <= 8'h38;
            13'h1DB8: rddata <= 8'h77;
            13'h1DB9: rddata <= 8'hCD;
            13'h1DBA: rddata <= 8'h1F;
            13'h1DBB: rddata <= 8'h1E;
            13'h1DBC: rddata <= 8'h18;
            13'h1DBD: rddata <= 8'h2C;
            13'h1DBE: rddata <= 8'hED;
            13'h1DBF: rddata <= 8'h5B;
            13'h1DC0: rddata <= 8'h00;
            13'h1DC1: rddata <= 8'h38;
            13'h1DC2: rddata <= 8'hAF;
            13'h1DC3: rddata <= 8'h57;
            13'h1DC4: rddata <= 8'hED;
            13'h1DC5: rddata <= 8'h52;
            13'h1DC6: rddata <= 8'h18;
            13'h1DC7: rddata <= 8'h1F;
            13'h1DC8: rddata <= 8'h11;
            13'h1DC9: rddata <= 8'hC0;
            13'h1DCA: rddata <= 8'h33;
            13'h1DCB: rddata <= 8'hE7;
            13'h1DCC: rddata <= 8'hD2;
            13'h1DCD: rddata <= 8'hD8;
            13'h1DCE: rddata <= 8'h1D;
            13'h1DCF: rddata <= 8'h11;
            13'h1DD0: rddata <= 8'h28;
            13'h1DD1: rddata <= 8'h00;
            13'h1DD2: rddata <= 8'h19;
            13'h1DD3: rddata <= 8'h22;
            13'h1DD4: rddata <= 8'h01;
            13'h1DD5: rddata <= 8'h38;
            13'h1DD6: rddata <= 8'h18;
            13'h1DD7: rddata <= 8'h12;
            13'h1DD8: rddata <= 8'hCD;
            13'h1DD9: rddata <= 8'hFE;
            13'h1DDA: rddata <= 8'h1D;
            13'h1DDB: rddata <= 8'h18;
            13'h1DDC: rddata <= 8'h0D;
            13'h1DDD: rddata <= 8'h3A;
            13'h1DDE: rddata <= 8'h00;
            13'h1DDF: rddata <= 8'h38;
            13'h1DE0: rddata <= 8'hB7;
            13'h1DE1: rddata <= 8'h28;
            13'h1DE2: rddata <= 8'h02;
            13'h1DE3: rddata <= 8'h2B;
            13'h1DE4: rddata <= 8'h3D;
            13'h1DE5: rddata <= 8'h36;
            13'h1DE6: rddata <= 8'h20;
            13'h1DE7: rddata <= 8'hCD;
            13'h1DE8: rddata <= 8'h3E;
            13'h1DE9: rddata <= 8'h1E;
            13'h1DEA: rddata <= 8'h2A;
            13'h1DEB: rddata <= 8'h01;
            13'h1DEC: rddata <= 8'h38;
            13'h1DED: rddata <= 8'h7E;
            13'h1DEE: rddata <= 8'h32;
            13'h1DEF: rddata <= 8'h0D;
            13'h1DF0: rddata <= 8'h38;
            13'h1DF1: rddata <= 8'h36;
            13'h1DF2: rddata <= 8'h7F;
            13'h1DF3: rddata <= 8'hD9;
            13'h1DF4: rddata <= 8'hF1;
            13'h1DF5: rddata <= 8'hC9;
            13'h1DF6: rddata <= 8'h2A;
            13'h1DF7: rddata <= 8'h01;
            13'h1DF8: rddata <= 8'h38;
            13'h1DF9: rddata <= 8'h3A;
            13'h1DFA: rddata <= 8'h0D;
            13'h1DFB: rddata <= 8'h38;
            13'h1DFC: rddata <= 8'h77;
            13'h1DFD: rddata <= 8'hC9;
            13'h1DFE: rddata <= 8'h01;
            13'h1DFF: rddata <= 8'h98;
            13'h1E00: rddata <= 8'h03;
            13'h1E01: rddata <= 8'h11;
            13'h1E02: rddata <= 8'h28;
            13'h1E03: rddata <= 8'h30;
            13'h1E04: rddata <= 8'h21;
            13'h1E05: rddata <= 8'h50;
            13'h1E06: rddata <= 8'h30;
            13'h1E07: rddata <= 8'hED;
            13'h1E08: rddata <= 8'hB0;
            13'h1E09: rddata <= 8'h06;
            13'h1E0A: rddata <= 8'h28;
            13'h1E0B: rddata <= 8'h21;
            13'h1E0C: rddata <= 8'hC1;
            13'h1E0D: rddata <= 8'h33;
            13'h1E0E: rddata <= 8'h36;
            13'h1E0F: rddata <= 8'h20;
            13'h1E10: rddata <= 8'h23;
            13'h1E11: rddata <= 8'h10;
            13'h1E12: rddata <= 8'hFB;
            13'h1E13: rddata <= 8'hC9;
            13'h1E14: rddata <= 8'h01;
            13'h1E15: rddata <= 8'hC8;
            13'h1E16: rddata <= 8'h00;
            13'h1E17: rddata <= 8'h11;
            13'h1E18: rddata <= 8'h32;
            13'h1E19: rddata <= 8'h00;
            13'h1E1A: rddata <= 8'hCD;
            13'h1E1B: rddata <= 8'h64;
            13'h1E1C: rddata <= 8'h1E;
            13'h1E1D: rddata <= 8'h18;
            13'h1E1E: rddata <= 8'hD4;
            13'h1E1F: rddata <= 8'h2A;
            13'h1E20: rddata <= 8'h01;
            13'h1E21: rddata <= 8'h38;
            13'h1E22: rddata <= 8'h3A;
            13'h1E23: rddata <= 8'h00;
            13'h1E24: rddata <= 8'h38;
            13'h1E25: rddata <= 8'h23;
            13'h1E26: rddata <= 8'h3C;
            13'h1E27: rddata <= 8'hFE;
            13'h1E28: rddata <= 8'h26;
            13'h1E29: rddata <= 8'h38;
            13'h1E2A: rddata <= 8'h13;
            13'h1E2B: rddata <= 8'h23;
            13'h1E2C: rddata <= 8'h23;
            13'h1E2D: rddata <= 8'h11;
            13'h1E2E: rddata <= 8'hE8;
            13'h1E2F: rddata <= 8'h33;
            13'h1E30: rddata <= 8'hE7;
            13'h1E31: rddata <= 8'h3E;
            13'h1E32: rddata <= 8'h00;
            13'h1E33: rddata <= 8'h38;
            13'h1E34: rddata <= 8'h09;
            13'h1E35: rddata <= 8'h21;
            13'h1E36: rddata <= 8'hC1;
            13'h1E37: rddata <= 8'h33;
            13'h1E38: rddata <= 8'hCD;
            13'h1E39: rddata <= 8'h3E;
            13'h1E3A: rddata <= 8'h1E;
            13'h1E3B: rddata <= 8'hC3;
            13'h1E3C: rddata <= 8'hFE;
            13'h1E3D: rddata <= 8'h1D;
            13'h1E3E: rddata <= 8'h22;
            13'h1E3F: rddata <= 8'h01;
            13'h1E40: rddata <= 8'h38;
            13'h1E41: rddata <= 8'h32;
            13'h1E42: rddata <= 8'h00;
            13'h1E43: rddata <= 8'h38;
            13'h1E44: rddata <= 8'hC9;
            13'h1E45: rddata <= 8'h06;
            13'h1E46: rddata <= 8'h20;
            13'h1E47: rddata <= 8'h21;
            13'h1E48: rddata <= 8'h00;
            13'h1E49: rddata <= 8'h30;
            13'h1E4A: rddata <= 8'hCD;
            13'h1E4B: rddata <= 8'h59;
            13'h1E4C: rddata <= 8'h1E;
            13'h1E4D: rddata <= 8'h06;
            13'h1E4E: rddata <= 8'h06;
            13'h1E4F: rddata <= 8'hCD;
            13'h1E50: rddata <= 8'h59;
            13'h1E51: rddata <= 8'h1E;
            13'h1E52: rddata <= 8'h21;
            13'h1E53: rddata <= 8'h29;
            13'h1E54: rddata <= 8'h30;
            13'h1E55: rddata <= 8'hAF;
            13'h1E56: rddata <= 8'hC3;
            13'h1E57: rddata <= 8'hE7;
            13'h1E58: rddata <= 8'h1D;
            13'h1E59: rddata <= 8'h11;
            13'h1E5A: rddata <= 8'hFF;
            13'h1E5B: rddata <= 8'h03;
            13'h1E5C: rddata <= 8'h70;
            13'h1E5D: rddata <= 8'h23;
            13'h1E5E: rddata <= 8'h1B;
            13'h1E5F: rddata <= 8'h7A;
            13'h1E60: rddata <= 8'hB3;
            13'h1E61: rddata <= 8'h20;
            13'h1E62: rddata <= 8'hF9;
            13'h1E63: rddata <= 8'hC9;
            13'h1E64: rddata <= 8'h78;
            13'h1E65: rddata <= 8'hB1;
            13'h1E66: rddata <= 8'hC8;
            13'h1E67: rddata <= 8'hAF;
            13'h1E68: rddata <= 8'hD3;
            13'h1E69: rddata <= 8'hFC;
            13'h1E6A: rddata <= 8'hCD;
            13'h1E6B: rddata <= 8'h76;
            13'h1E6C: rddata <= 8'h1E;
            13'h1E6D: rddata <= 8'h3C;
            13'h1E6E: rddata <= 8'hD3;
            13'h1E6F: rddata <= 8'hFC;
            13'h1E70: rddata <= 8'hCD;
            13'h1E71: rddata <= 8'h76;
            13'h1E72: rddata <= 8'h1E;
            13'h1E73: rddata <= 8'h0B;
            13'h1E74: rddata <= 8'h18;
            13'h1E75: rddata <= 8'hEE;
            13'h1E76: rddata <= 8'hD5;
            13'h1E77: rddata <= 8'hE1;
            13'h1E78: rddata <= 8'h7C;
            13'h1E79: rddata <= 8'hB5;
            13'h1E7A: rddata <= 8'hC8;
            13'h1E7B: rddata <= 8'h2B;
            13'h1E7C: rddata <= 8'h18;
            13'h1E7D: rddata <= 8'hFA;
            13'h1E7E: rddata <= 8'hF7;
            13'h1E7F: rddata <= 8'h12;
            13'h1E80: rddata <= 8'hD9;
            13'h1E81: rddata <= 8'h2A;
            13'h1E82: rddata <= 8'h0B;
            13'h1E83: rddata <= 8'h38;
            13'h1E84: rddata <= 8'h7C;
            13'h1E85: rddata <= 8'hB7;
            13'h1E86: rddata <= 8'h28;
            13'h1E87: rddata <= 8'h1A;
            13'h1E88: rddata <= 8'hEB;
            13'h1E89: rddata <= 8'h21;
            13'h1E8A: rddata <= 8'h0F;
            13'h1E8B: rddata <= 8'h38;
            13'h1E8C: rddata <= 8'h34;
            13'h1E8D: rddata <= 8'h7E;
            13'h1E8E: rddata <= 8'hFE;
            13'h1E8F: rddata <= 8'h0F;
            13'h1E90: rddata <= 8'h38;
            13'h1E91: rddata <= 8'h3C;
            13'h1E92: rddata <= 8'h36;
            13'h1E93: rddata <= 8'h05;
            13'h1E94: rddata <= 8'hEB;
            13'h1E95: rddata <= 8'h23;
            13'h1E96: rddata <= 8'h7E;
            13'h1E97: rddata <= 8'h22;
            13'h1E98: rddata <= 8'h0B;
            13'h1E99: rddata <= 8'h38;
            13'h1E9A: rddata <= 8'hB7;
            13'h1E9B: rddata <= 8'hF2;
            13'h1E9C: rddata <= 8'h36;
            13'h1E9D: rddata <= 8'h1F;
            13'h1E9E: rddata <= 8'hAF;
            13'h1E9F: rddata <= 8'h32;
            13'h1EA0: rddata <= 8'h0C;
            13'h1EA1: rddata <= 8'h38;
            13'h1EA2: rddata <= 8'h01;
            13'h1EA3: rddata <= 8'hFF;
            13'h1EA4: rddata <= 8'h00;
            13'h1EA5: rddata <= 8'hED;
            13'h1EA6: rddata <= 8'h78;
            13'h1EA7: rddata <= 8'h2F;
            13'h1EA8: rddata <= 8'hE6;
            13'h1EA9: rddata <= 8'h3F;
            13'h1EAA: rddata <= 8'h21;
            13'h1EAB: rddata <= 8'h0E;
            13'h1EAC: rddata <= 8'h38;
            13'h1EAD: rddata <= 8'h28;
            13'h1EAE: rddata <= 8'h16;
            13'h1EAF: rddata <= 8'h06;
            13'h1EB0: rddata <= 8'h7F;
            13'h1EB1: rddata <= 8'hED;
            13'h1EB2: rddata <= 8'h78;
            13'h1EB3: rddata <= 8'h2F;
            13'h1EB4: rddata <= 8'hE6;
            13'h1EB5: rddata <= 8'h0F;
            13'h1EB6: rddata <= 8'h20;
            13'h1EB7: rddata <= 8'h1F;
            13'h1EB8: rddata <= 8'h06;
            13'h1EB9: rddata <= 8'hBF;
            13'h1EBA: rddata <= 8'hED;
            13'h1EBB: rddata <= 8'h78;
            13'h1EBC: rddata <= 8'h2F;
            13'h1EBD: rddata <= 8'hE6;
            13'h1EBE: rddata <= 8'h3F;
            13'h1EBF: rddata <= 8'h20;
            13'h1EC0: rddata <= 8'h16;
            13'h1EC1: rddata <= 8'hCB;
            13'h1EC2: rddata <= 8'h08;
            13'h1EC3: rddata <= 8'h38;
            13'h1EC4: rddata <= 8'hF5;
            13'h1EC5: rddata <= 8'h23;
            13'h1EC6: rddata <= 8'h3E;
            13'h1EC7: rddata <= 8'h46;
            13'h1EC8: rddata <= 8'hBE;
            13'h1EC9: rddata <= 8'h38;
            13'h1ECA: rddata <= 8'h03;
            13'h1ECB: rddata <= 8'h28;
            13'h1ECC: rddata <= 8'h04;
            13'h1ECD: rddata <= 8'h34;
            13'h1ECE: rddata <= 8'hAF;
            13'h1ECF: rddata <= 8'hD9;
            13'h1ED0: rddata <= 8'hC9;
            13'h1ED1: rddata <= 8'h34;
            13'h1ED2: rddata <= 8'h2B;
            13'h1ED3: rddata <= 8'h36;
            13'h1ED4: rddata <= 8'h00;
            13'h1ED5: rddata <= 8'h18;
            13'h1ED6: rddata <= 8'hF7;
            13'h1ED7: rddata <= 8'h11;
            13'h1ED8: rddata <= 8'h00;
            13'h1ED9: rddata <= 8'h00;
            13'h1EDA: rddata <= 8'h1C;
            13'h1EDB: rddata <= 8'h1F;
            13'h1EDC: rddata <= 8'h30;
            13'h1EDD: rddata <= 8'hFC;
            13'h1EDE: rddata <= 8'h7B;
            13'h1EDF: rddata <= 8'hCB;
            13'h1EE0: rddata <= 8'h18;
            13'h1EE1: rddata <= 8'h30;
            13'h1EE2: rddata <= 8'h04;
            13'h1EE3: rddata <= 8'hC6;
            13'h1EE4: rddata <= 8'h06;
            13'h1EE5: rddata <= 8'h18;
            13'h1EE6: rddata <= 8'hF8;
            13'h1EE7: rddata <= 8'h5F;
            13'h1EE8: rddata <= 8'hBE;
            13'h1EE9: rddata <= 8'h77;
            13'h1EEA: rddata <= 8'h23;
            13'h1EEB: rddata <= 8'h20;
            13'h1EEC: rddata <= 8'h0F;
            13'h1EED: rddata <= 8'h3E;
            13'h1EEE: rddata <= 8'h04;
            13'h1EEF: rddata <= 8'hBE;
            13'h1EF0: rddata <= 8'h38;
            13'h1EF1: rddata <= 8'h05;
            13'h1EF2: rddata <= 8'h28;
            13'h1EF3: rddata <= 8'h0C;
            13'h1EF4: rddata <= 8'h34;
            13'h1EF5: rddata <= 8'h18;
            13'h1EF6: rddata <= 8'h02;
            13'h1EF7: rddata <= 8'h36;
            13'h1EF8: rddata <= 8'h06;
            13'h1EF9: rddata <= 8'hAF;
            13'h1EFA: rddata <= 8'hD9;
            13'h1EFB: rddata <= 8'hC9;
            13'h1EFC: rddata <= 8'h36;
            13'h1EFD: rddata <= 8'h00;
            13'h1EFE: rddata <= 8'h18;
            13'h1EFF: rddata <= 8'hF9;
            13'h1F00: rddata <= 8'h34;
            13'h1F01: rddata <= 8'h06;
            13'h1F02: rddata <= 8'h7F;
            13'h1F03: rddata <= 8'hED;
            13'h1F04: rddata <= 8'h78;
            13'h1F05: rddata <= 8'hCB;
            13'h1F06: rddata <= 8'h6F;
            13'h1F07: rddata <= 8'hDD;
            13'h1F08: rddata <= 8'h21;
            13'h1F09: rddata <= 8'h93;
            13'h1F0A: rddata <= 8'h1F;
            13'h1F0B: rddata <= 8'h28;
            13'h1F0C: rddata <= 8'h0C;
            13'h1F0D: rddata <= 8'hCB;
            13'h1F0E: rddata <= 8'h67;
            13'h1F0F: rddata <= 8'hDD;
            13'h1F10: rddata <= 8'h21;
            13'h1F11: rddata <= 8'h65;
            13'h1F12: rddata <= 8'h1F;
            13'h1F13: rddata <= 8'h28;
            13'h1F14: rddata <= 8'h04;
            13'h1F15: rddata <= 8'hDD;
            13'h1F16: rddata <= 8'h21;
            13'h1F17: rddata <= 8'h37;
            13'h1F18: rddata <= 8'h1F;
            13'h1F19: rddata <= 8'hDD;
            13'h1F1A: rddata <= 8'h19;
            13'h1F1B: rddata <= 8'hDD;
            13'h1F1C: rddata <= 8'h7E;
            13'h1F1D: rddata <= 8'h00;
            13'h1F1E: rddata <= 8'hB7;
            13'h1F1F: rddata <= 8'hF2;
            13'h1F20: rddata <= 8'h36;
            13'h1F21: rddata <= 8'h1F;
            13'h1F22: rddata <= 8'hD6;
            13'h1F23: rddata <= 8'h7F;
            13'h1F24: rddata <= 8'h4F;
            13'h1F25: rddata <= 8'h21;
            13'h1F26: rddata <= 8'h44;
            13'h1F27: rddata <= 8'h02;
            13'h1F28: rddata <= 8'h23;
            13'h1F29: rddata <= 8'h7E;
            13'h1F2A: rddata <= 8'hB7;
            13'h1F2B: rddata <= 8'hF2;
            13'h1F2C: rddata <= 8'h28;
            13'h1F2D: rddata <= 8'h1F;
            13'h1F2E: rddata <= 8'h0D;
            13'h1F2F: rddata <= 8'h20;
            13'h1F30: rddata <= 8'hF7;
            13'h1F31: rddata <= 8'h22;
            13'h1F32: rddata <= 8'h0B;
            13'h1F33: rddata <= 8'h38;
            13'h1F34: rddata <= 8'hE6;
            13'h1F35: rddata <= 8'h7F;
            13'h1F36: rddata <= 8'hD9;
            13'h1F37: rddata <= 8'hC9;
            13'h1F38: rddata <= 8'h3D;
            13'h1F39: rddata <= 8'h08;
            13'h1F3A: rddata <= 8'h3A;
            13'h1F3B: rddata <= 8'h0D;
            13'h1F3C: rddata <= 8'h3B;
            13'h1F3D: rddata <= 8'h2E;
            13'h1F3E: rddata <= 8'h2D;
            13'h1F3F: rddata <= 8'h2F;
            13'h1F40: rddata <= 8'h30;
            13'h1F41: rddata <= 8'h70;
            13'h1F42: rddata <= 8'h6C;
            13'h1F43: rddata <= 8'h2C;
            13'h1F44: rddata <= 8'h39;
            13'h1F45: rddata <= 8'h6F;
            13'h1F46: rddata <= 8'h6B;
            13'h1F47: rddata <= 8'h6D;
            13'h1F48: rddata <= 8'h6E;
            13'h1F49: rddata <= 8'h6A;
            13'h1F4A: rddata <= 8'h38;
            13'h1F4B: rddata <= 8'h69;
            13'h1F4C: rddata <= 8'h37;
            13'h1F4D: rddata <= 8'h75;
            13'h1F4E: rddata <= 8'h68;
            13'h1F4F: rddata <= 8'h62;
            13'h1F50: rddata <= 8'h36;
            13'h1F51: rddata <= 8'h79;
            13'h1F52: rddata <= 8'h67;
            13'h1F53: rddata <= 8'h76;
            13'h1F54: rddata <= 8'h63;
            13'h1F55: rddata <= 8'h66;
            13'h1F56: rddata <= 8'h35;
            13'h1F57: rddata <= 8'h74;
            13'h1F58: rddata <= 8'h34;
            13'h1F59: rddata <= 8'h72;
            13'h1F5A: rddata <= 8'h64;
            13'h1F5B: rddata <= 8'h78;
            13'h1F5C: rddata <= 8'h33;
            13'h1F5D: rddata <= 8'h65;
            13'h1F5E: rddata <= 8'h73;
            13'h1F5F: rddata <= 8'h7A;
            13'h1F60: rddata <= 8'h20;
            13'h1F61: rddata <= 8'h61;
            13'h1F62: rddata <= 8'h32;
            13'h1F63: rddata <= 8'h77;
            13'h1F64: rddata <= 8'h31;
            13'h1F65: rddata <= 8'h71;
            13'h1F66: rddata <= 8'h2B;
            13'h1F67: rddata <= 8'h5C;
            13'h1F68: rddata <= 8'h2A;
            13'h1F69: rddata <= 8'h0D;
            13'h1F6A: rddata <= 8'h40;
            13'h1F6B: rddata <= 8'h3E;
            13'h1F6C: rddata <= 8'h5F;
            13'h1F6D: rddata <= 8'h5E;
            13'h1F6E: rddata <= 8'h3F;
            13'h1F6F: rddata <= 8'h50;
            13'h1F70: rddata <= 8'h4C;
            13'h1F71: rddata <= 8'h3C;
            13'h1F72: rddata <= 8'h29;
            13'h1F73: rddata <= 8'h4F;
            13'h1F74: rddata <= 8'h4B;
            13'h1F75: rddata <= 8'h4D;
            13'h1F76: rddata <= 8'h4E;
            13'h1F77: rddata <= 8'h4A;
            13'h1F78: rddata <= 8'h28;
            13'h1F79: rddata <= 8'h49;
            13'h1F7A: rddata <= 8'h27;
            13'h1F7B: rddata <= 8'h55;
            13'h1F7C: rddata <= 8'h48;
            13'h1F7D: rddata <= 8'h42;
            13'h1F7E: rddata <= 8'h26;
            13'h1F7F: rddata <= 8'h59;
            13'h1F80: rddata <= 8'h47;
            13'h1F81: rddata <= 8'h56;
            13'h1F82: rddata <= 8'h43;
            13'h1F83: rddata <= 8'h46;
            13'h1F84: rddata <= 8'h25;
            13'h1F85: rddata <= 8'h54;
            13'h1F86: rddata <= 8'h24;
            13'h1F87: rddata <= 8'h52;
            13'h1F88: rddata <= 8'h44;
            13'h1F89: rddata <= 8'h58;
            13'h1F8A: rddata <= 8'h23;
            13'h1F8B: rddata <= 8'h45;
            13'h1F8C: rddata <= 8'h53;
            13'h1F8D: rddata <= 8'h5A;
            13'h1F8E: rddata <= 8'h20;
            13'h1F8F: rddata <= 8'h41;
            13'h1F90: rddata <= 8'h22;
            13'h1F91: rddata <= 8'h57;
            13'h1F92: rddata <= 8'h21;
            13'h1F93: rddata <= 8'h51;
            13'h1F94: rddata <= 8'h82;
            13'h1F95: rddata <= 8'h1C;
            13'h1F96: rddata <= 8'hC1;
            13'h1F97: rddata <= 8'h0D;
            13'h1F98: rddata <= 8'h94;
            13'h1F99: rddata <= 8'hC4;
            13'h1F9A: rddata <= 8'h81;
            13'h1F9B: rddata <= 8'h1E;
            13'h1F9C: rddata <= 8'h30;
            13'h1F9D: rddata <= 8'h10;
            13'h1F9E: rddata <= 8'hCA;
            13'h1F9F: rddata <= 8'hC3;
            13'h1FA0: rddata <= 8'h92;
            13'h1FA1: rddata <= 8'h0F;
            13'h1FA2: rddata <= 8'h9D;
            13'h1FA3: rddata <= 8'h0D;
            13'h1FA4: rddata <= 8'hC8;
            13'h1FA5: rddata <= 8'h9C;
            13'h1FA6: rddata <= 8'h8D;
            13'h1FA7: rddata <= 8'h09;
            13'h1FA8: rddata <= 8'h8C;
            13'h1FA9: rddata <= 8'h15;
            13'h1FAA: rddata <= 8'h08;
            13'h1FAB: rddata <= 8'hC9;
            13'h1FAC: rddata <= 8'h90;
            13'h1FAD: rddata <= 8'h19;
            13'h1FAE: rddata <= 8'h07;
            13'h1FAF: rddata <= 8'hC7;
            13'h1FB0: rddata <= 8'h03;
            13'h1FB1: rddata <= 8'h83;
            13'h1FB2: rddata <= 8'h88;
            13'h1FB3: rddata <= 8'h84;
            13'h1FB4: rddata <= 8'hA5;
            13'h1FB5: rddata <= 8'h12;
            13'h1FB6: rddata <= 8'h86;
            13'h1FB7: rddata <= 8'h18;
            13'h1FB8: rddata <= 8'h8A;
            13'h1FB9: rddata <= 8'h85;
            13'h1FBA: rddata <= 8'h13;
            13'h1FBB: rddata <= 8'h9A;
            13'h1FBC: rddata <= 8'hC6;
            13'h1FBD: rddata <= 8'h9B;
            13'h1FBE: rddata <= 8'h97;
            13'h1FBF: rddata <= 8'h8E;
            13'h1FC0: rddata <= 8'h89;
            13'h1FC1: rddata <= 8'h11;
            13'h1FC2: rddata <= 8'hE5;
            13'h1FC3: rddata <= 8'h21;
            13'h1FC4: rddata <= 8'h04;
            13'h1FC5: rddata <= 8'h00;
            13'h1FC6: rddata <= 8'h39;
            13'h1FC7: rddata <= 8'h22;
            13'h1FC8: rddata <= 8'hF9;
            13'h1FC9: rddata <= 8'h38;
            13'h1FCA: rddata <= 8'hE1;
            13'h1FCB: rddata <= 8'hC3;
            13'h1FCC: rddata <= 8'h25;
            13'h1FCD: rddata <= 8'h1A;
            13'h1FCE: rddata <= 8'h2A;
            13'h1FCF: rddata <= 8'hF9;
            13'h1FD0: rddata <= 8'h38;
            13'h1FD1: rddata <= 8'hF9;
            13'h1FD2: rddata <= 8'h2A;
            13'h1FD3: rddata <= 8'hCE;
            13'h1FD4: rddata <= 8'h38;
            13'h1FD5: rddata <= 8'hCD;
            13'h1FD6: rddata <= 8'h20;
            13'h1FD7: rddata <= 8'h0C;
            13'h1FD8: rddata <= 8'h2B;
            13'h1FD9: rddata <= 8'h2B;
            13'h1FDA: rddata <= 8'h22;
            13'h1FDB: rddata <= 8'hF9;
            13'h1FDC: rddata <= 8'h38;
            13'h1FDD: rddata <= 8'h21;
            13'h1FDE: rddata <= 8'hB1;
            13'h1FDF: rddata <= 8'h38;
            13'h1FE0: rddata <= 8'hC9;
            13'h1FE1: rddata <= 8'h3E;
            13'h1FE2: rddata <= 8'hFF;
            13'h1FE3: rddata <= 8'hD3;
            13'h1FE4: rddata <= 8'hFE;
            13'h1FE5: rddata <= 8'hC3;
            13'h1FE6: rddata <= 8'h41;
            13'h1FE7: rddata <= 8'h00;
            13'h1FE8: rddata <= 8'h3E;
            13'h1FE9: rddata <= 8'hAA;
            13'h1FEA: rddata <= 8'hD3;
            13'h1FEB: rddata <= 8'hFF;
            13'h1FEC: rddata <= 8'h32;
            13'h1FED: rddata <= 8'h09;
            13'h1FEE: rddata <= 8'h38;
            13'h1FEF: rddata <= 8'hC3;
            13'h1FF0: rddata <= 8'h10;
            13'h1FF1: rddata <= 8'h20;
            13'h1FF2: rddata <= 8'h21;
            13'h1FF3: rddata <= 8'h5F;
            13'h1FF4: rddata <= 8'h01;
            13'h1FF5: rddata <= 8'hC3;
            13'h1FF6: rddata <= 8'h9D;
            13'h1FF7: rddata <= 8'h0E;
            13'h1FF8: rddata <= 8'hF5;
            13'h1FF9: rddata <= 8'hF5;
            13'h1FFA: rddata <= 8'hF5;
            13'h1FFB: rddata <= 8'hF5;
            13'h1FFC: rddata <= 8'hF5;
            13'h1FFD: rddata <= 8'hF5;
            13'h1FFE: rddata <= 8'hF5;
            13'h1FFF: rddata <= 8'hF5;
            default:  rddata <= 8'h00; // NOP
        endcase

endmodule
